`timescale 1ns / 1ps

//数据存储器，是RAM，有写入功能


module data_mem( 
    input [9:0] addr,//需要访问的地址（10位）
    input [3:0] led_addr,
    input [31:0] din,//数据
    input [3:0] mode, //sel
    input clk,//时钟输入端
    input WE,//存储：当为1时从存储端输入数据
    input clr,//清空：当为1时，重置内存为0
    output [31:0] dout,//从地址加载的数据（32位）
    output [31:0] led_data_out
);

// module RAM( addr,led_addr ,din,mode,clk , WE,,clr,dout , led_data_out);
// input [9:0] addr;
// input [3:0] led_addr,
// input [31:0] din;
// input [3:0] mode;
// input WE,clk,clr;
// output [31:0] dout;
// output [31:0] led_data_out
//?20 位地址？？这里实现的是10位地址
reg [7:0] mem1[1023:0], mem2[1023:0],mem3[1023:0],mem4[1023:0];
// reg  [31:0] dout;



assign dout = {
    mem4[addr], 
    mem3[addr],
    mem2[addr],
    mem1[addr]
};
assign  led_data_out = {
    mem4[led_addr], 
    mem3[led_addr],
    mem2[led_addr],
    mem1[led_addr]
}

// }{[7:0] <= 
//     dout[15:8] <= 
//     dout[23:16] <= 
//     dout[31:24] <= ;

always@(posedge clk )
begin

if(WE)
  begin
        // mem1[addr[21:2]] <= din[7:0];
        //   mem2[addr[21:2]] <= din[15:8];
        //   mem3[addr[21:2]] <= din[23:16];
        //   mem4[addr[21:2]] <= din[31:24];

    case(mode)
    4'b1111:
    begin
        mem1[addr] <= din[7:0];
        mem2[addr] <= din[15:8];
        mem3[addr] <= din[23:16];
        mem4[addr] <= din[31:24];
    end
    4'b0001:
    begin
        mem1[addr] <= din[7:0];
    end
    4'b0010:
    begin
        mem2[addr] <= din[15:8];
    end
    4'b0100:
    begin
        mem3[addr] <= din[23:16];
    end
    4'b1000:
    begin
        mem4[addr] <= din[31:24];
    end
    4'b0011:
    begin
        mem1[addr] <= din[7:0];
        mem2[addr] <= din[15:8];    
    end
    4'b1100:
    begin
        mem3[addr] <= din[23:16];
        mem4[addr] <= din[31:24];
    end

  end
end  




initial
begin
mem1[0]<=0;  mem2[0]<=0; mem3[0]<=0; mem4[0]<=0;
mem1[1]<=0;  mem2[1]<=0; mem3[1]<=0; mem4[1]<=0;
mem1[2]<=0;  mem2[2]<=0; mem3[2]<=0; mem4[2]<=0;
mem1[3]<=0;  mem2[3]<=0; mem3[3]<=0; mem4[3]<=0;
mem1[4]<=0;  mem2[4]<=0; mem3[4]<=0; mem4[4]<=0;
mem1[5]<=0;  mem2[5]<=0; mem3[5]<=0; mem4[5]<=0;
mem1[6]<=0;  mem2[6]<=0; mem3[6]<=0; mem4[6]<=0;
mem1[7]<=0;  mem2[7]<=0; mem3[7]<=0; mem4[7]<=0;
mem1[8]<=0;  mem2[8]<=0; mem3[8]<=0; mem4[8]<=0;
mem1[9]<=0;  mem2[9]<=0; mem3[9]<=0; mem4[9]<=0;
mem1[10]<=0;  mem2[10]<=0; mem3[10]<=0; mem4[10]<=0;
mem1[11]<=0;  mem2[11]<=0; mem3[11]<=0; mem4[11]<=0;
mem1[12]<=0;  mem2[12]<=0; mem3[12]<=0; mem4[12]<=0;
mem1[13]<=0;  mem2[13]<=0; mem3[13]<=0; mem4[13]<=0;
mem1[14]<=0;  mem2[14]<=0; mem3[14]<=0; mem4[14]<=0;
mem1[15]<=0;  mem2[15]<=0; mem3[15]<=0; mem4[15]<=0;
mem1[16]<=0;  mem2[16]<=0; mem3[16]<=0; mem4[16]<=0;
mem1[17]<=0;  mem2[17]<=0; mem3[17]<=0; mem4[17]<=0;
mem1[18]<=0;  mem2[18]<=0; mem3[18]<=0; mem4[18]<=0;
mem1[19]<=0;  mem2[19]<=0; mem3[19]<=0; mem4[19]<=0;
mem1[20]<=0;  mem2[20]<=0; mem3[20]<=0; mem4[20]<=0;
mem1[21]<=0;  mem2[21]<=0; mem3[21]<=0; mem4[21]<=0;
mem1[22]<=0;  mem2[22]<=0; mem3[22]<=0; mem4[22]<=0;
mem1[23]<=0;  mem2[23]<=0; mem3[23]<=0; mem4[23]<=0;
mem1[24]<=0;  mem2[24]<=0; mem3[24]<=0; mem4[24]<=0;
mem1[25]<=0;  mem2[25]<=0; mem3[25]<=0; mem4[25]<=0;
mem1[26]<=0;  mem2[26]<=0; mem3[26]<=0; mem4[26]<=0;
mem1[27]<=0;  mem2[27]<=0; mem3[27]<=0; mem4[27]<=0;
mem1[28]<=0;  mem2[28]<=0; mem3[28]<=0; mem4[28]<=0;
mem1[29]<=0;  mem2[29]<=0; mem3[29]<=0; mem4[29]<=0;
mem1[30]<=0;  mem2[30]<=0; mem3[30]<=0; mem4[30]<=0;
mem1[31]<=0;  mem2[31]<=0; mem3[31]<=0; mem4[31]<=0;
mem1[32]<=0;  mem2[32]<=0; mem3[32]<=0; mem4[32]<=0;
mem1[33]<=0;  mem2[33]<=0; mem3[33]<=0; mem4[33]<=0;
mem1[34]<=0;  mem2[34]<=0; mem3[34]<=0; mem4[34]<=0;
mem1[35]<=0;  mem2[35]<=0; mem3[35]<=0; mem4[35]<=0;
mem1[36]<=0;  mem2[36]<=0; mem3[36]<=0; mem4[36]<=0;
mem1[37]<=0;  mem2[37]<=0; mem3[37]<=0; mem4[37]<=0;
mem1[38]<=0;  mem2[38]<=0; mem3[38]<=0; mem4[38]<=0;
mem1[39]<=0;  mem2[39]<=0; mem3[39]<=0; mem4[39]<=0;
mem1[40]<=0;  mem2[40]<=0; mem3[40]<=0; mem4[40]<=0;
mem1[41]<=0;  mem2[41]<=0; mem3[41]<=0; mem4[41]<=0;
mem1[42]<=0;  mem2[42]<=0; mem3[42]<=0; mem4[42]<=0;
mem1[43]<=0;  mem2[43]<=0; mem3[43]<=0; mem4[43]<=0;
mem1[44]<=0;  mem2[44]<=0; mem3[44]<=0; mem4[44]<=0;
mem1[45]<=0;  mem2[45]<=0; mem3[45]<=0; mem4[45]<=0;
mem1[46]<=0;  mem2[46]<=0; mem3[46]<=0; mem4[46]<=0;
mem1[47]<=0;  mem2[47]<=0; mem3[47]<=0; mem4[47]<=0;
mem1[48]<=0;  mem2[48]<=0; mem3[48]<=0; mem4[48]<=0;
mem1[49]<=0;  mem2[49]<=0; mem3[49]<=0; mem4[49]<=0;
mem1[50]<=0;  mem2[50]<=0; mem3[50]<=0; mem4[50]<=0;
mem1[51]<=0;  mem2[51]<=0; mem3[51]<=0; mem4[51]<=0;
mem1[52]<=0;  mem2[52]<=0; mem3[52]<=0; mem4[52]<=0;
mem1[53]<=0;  mem2[53]<=0; mem3[53]<=0; mem4[53]<=0;
mem1[54]<=0;  mem2[54]<=0; mem3[54]<=0; mem4[54]<=0;
mem1[55]<=0;  mem2[55]<=0; mem3[55]<=0; mem4[55]<=0;
mem1[56]<=0;  mem2[56]<=0; mem3[56]<=0; mem4[56]<=0;
mem1[57]<=0;  mem2[57]<=0; mem3[57]<=0; mem4[57]<=0;
mem1[58]<=0;  mem2[58]<=0; mem3[58]<=0; mem4[58]<=0;
mem1[59]<=0;  mem2[59]<=0; mem3[59]<=0; mem4[59]<=0;
mem1[60]<=0;  mem2[60]<=0; mem3[60]<=0; mem4[60]<=0;
mem1[61]<=0;  mem2[61]<=0; mem3[61]<=0; mem4[61]<=0;
mem1[62]<=0;  mem2[62]<=0; mem3[62]<=0; mem4[62]<=0;
mem1[63]<=0;  mem2[63]<=0; mem3[63]<=0; mem4[63]<=0;
mem1[64]<=0;  mem2[64]<=0; mem3[64]<=0; mem4[64]<=0;
mem1[65]<=0;  mem2[65]<=0; mem3[65]<=0; mem4[65]<=0;
mem1[66]<=0;  mem2[66]<=0; mem3[66]<=0; mem4[66]<=0;
mem1[67]<=0;  mem2[67]<=0; mem3[67]<=0; mem4[67]<=0;
mem1[68]<=0;  mem2[68]<=0; mem3[68]<=0; mem4[68]<=0;
mem1[69]<=0;  mem2[69]<=0; mem3[69]<=0; mem4[69]<=0;
mem1[70]<=0;  mem2[70]<=0; mem3[70]<=0; mem4[70]<=0;
mem1[71]<=0;  mem2[71]<=0; mem3[71]<=0; mem4[71]<=0;
mem1[72]<=0;  mem2[72]<=0; mem3[72]<=0; mem4[72]<=0;
mem1[73]<=0;  mem2[73]<=0; mem3[73]<=0; mem4[73]<=0;
mem1[74]<=0;  mem2[74]<=0; mem3[74]<=0; mem4[74]<=0;
mem1[75]<=0;  mem2[75]<=0; mem3[75]<=0; mem4[75]<=0;
mem1[76]<=0;  mem2[76]<=0; mem3[76]<=0; mem4[76]<=0;
mem1[77]<=0;  mem2[77]<=0; mem3[77]<=0; mem4[77]<=0;
mem1[78]<=0;  mem2[78]<=0; mem3[78]<=0; mem4[78]<=0;
mem1[79]<=0;  mem2[79]<=0; mem3[79]<=0; mem4[79]<=0;
mem1[80]<=0;  mem2[80]<=0; mem3[80]<=0; mem4[80]<=0;
mem1[81]<=0;  mem2[81]<=0; mem3[81]<=0; mem4[81]<=0;
mem1[82]<=0;  mem2[82]<=0; mem3[82]<=0; mem4[82]<=0;
mem1[83]<=0;  mem2[83]<=0; mem3[83]<=0; mem4[83]<=0;
mem1[84]<=0;  mem2[84]<=0; mem3[84]<=0; mem4[84]<=0;
mem1[85]<=0;  mem2[85]<=0; mem3[85]<=0; mem4[85]<=0;
mem1[86]<=0;  mem2[86]<=0; mem3[86]<=0; mem4[86]<=0;
mem1[87]<=0;  mem2[87]<=0; mem3[87]<=0; mem4[87]<=0;
mem1[88]<=0;  mem2[88]<=0; mem3[88]<=0; mem4[88]<=0;
mem1[89]<=0;  mem2[89]<=0; mem3[89]<=0; mem4[89]<=0;
mem1[90]<=0;  mem2[90]<=0; mem3[90]<=0; mem4[90]<=0;
mem1[91]<=0;  mem2[91]<=0; mem3[91]<=0; mem4[91]<=0;
mem1[92]<=0;  mem2[92]<=0; mem3[92]<=0; mem4[92]<=0;
mem1[93]<=0;  mem2[93]<=0; mem3[93]<=0; mem4[93]<=0;
mem1[94]<=0;  mem2[94]<=0; mem3[94]<=0; mem4[94]<=0;
mem1[95]<=0;  mem2[95]<=0; mem3[95]<=0; mem4[95]<=0;
mem1[96]<=0;  mem2[96]<=0; mem3[96]<=0; mem4[96]<=0;
mem1[97]<=0;  mem2[97]<=0; mem3[97]<=0; mem4[97]<=0;
mem1[98]<=0;  mem2[98]<=0; mem3[98]<=0; mem4[98]<=0;
mem1[99]<=0;  mem2[99]<=0; mem3[99]<=0; mem4[99]<=0;
mem1[100]<=0;  mem2[100]<=0; mem3[100]<=0; mem4[100]<=0;
mem1[101]<=0;  mem2[101]<=0; mem3[101]<=0; mem4[101]<=0;
mem1[102]<=0;  mem2[102]<=0; mem3[102]<=0; mem4[102]<=0;
mem1[103]<=0;  mem2[103]<=0; mem3[103]<=0; mem4[103]<=0;
mem1[104]<=0;  mem2[104]<=0; mem3[104]<=0; mem4[104]<=0;
mem1[105]<=0;  mem2[105]<=0; mem3[105]<=0; mem4[105]<=0;
mem1[106]<=0;  mem2[106]<=0; mem3[106]<=0; mem4[106]<=0;
mem1[107]<=0;  mem2[107]<=0; mem3[107]<=0; mem4[107]<=0;
mem1[108]<=0;  mem2[108]<=0; mem3[108]<=0; mem4[108]<=0;
mem1[109]<=0;  mem2[109]<=0; mem3[109]<=0; mem4[109]<=0;
mem1[110]<=0;  mem2[110]<=0; mem3[110]<=0; mem4[110]<=0;
mem1[111]<=0;  mem2[111]<=0; mem3[111]<=0; mem4[111]<=0;
mem1[112]<=0;  mem2[112]<=0; mem3[112]<=0; mem4[112]<=0;
mem1[113]<=0;  mem2[113]<=0; mem3[113]<=0; mem4[113]<=0;
mem1[114]<=0;  mem2[114]<=0; mem3[114]<=0; mem4[114]<=0;
mem1[115]<=0;  mem2[115]<=0; mem3[115]<=0; mem4[115]<=0;
mem1[116]<=0;  mem2[116]<=0; mem3[116]<=0; mem4[116]<=0;
mem1[117]<=0;  mem2[117]<=0; mem3[117]<=0; mem4[117]<=0;
mem1[118]<=0;  mem2[118]<=0; mem3[118]<=0; mem4[118]<=0;
mem1[119]<=0;  mem2[119]<=0; mem3[119]<=0; mem4[119]<=0;
mem1[120]<=0;  mem2[120]<=0; mem3[120]<=0; mem4[120]<=0;
mem1[121]<=0;  mem2[121]<=0; mem3[121]<=0; mem4[121]<=0;
mem1[122]<=0;  mem2[122]<=0; mem3[122]<=0; mem4[122]<=0;
mem1[123]<=0;  mem2[123]<=0; mem3[123]<=0; mem4[123]<=0;
mem1[124]<=0;  mem2[124]<=0; mem3[124]<=0; mem4[124]<=0;
mem1[125]<=0;  mem2[125]<=0; mem3[125]<=0; mem4[125]<=0;
mem1[126]<=0;  mem2[126]<=0; mem3[126]<=0; mem4[126]<=0;
mem1[127]<=0;  mem2[127]<=0; mem3[127]<=0; mem4[127]<=0;
mem1[128]<=0;  mem2[128]<=0; mem3[128]<=0; mem4[128]<=0;
mem1[129]<=0;  mem2[129]<=0; mem3[129]<=0; mem4[129]<=0;
mem1[130]<=0;  mem2[130]<=0; mem3[130]<=0; mem4[130]<=0;
mem1[131]<=0;  mem2[131]<=0; mem3[131]<=0; mem4[131]<=0;
mem1[132]<=0;  mem2[132]<=0; mem3[132]<=0; mem4[132]<=0;
mem1[133]<=0;  mem2[133]<=0; mem3[133]<=0; mem4[133]<=0;
mem1[134]<=0;  mem2[134]<=0; mem3[134]<=0; mem4[134]<=0;
mem1[135]<=0;  mem2[135]<=0; mem3[135]<=0; mem4[135]<=0;
mem1[136]<=0;  mem2[136]<=0; mem3[136]<=0; mem4[136]<=0;
mem1[137]<=0;  mem2[137]<=0; mem3[137]<=0; mem4[137]<=0;
mem1[138]<=0;  mem2[138]<=0; mem3[138]<=0; mem4[138]<=0;
mem1[139]<=0;  mem2[139]<=0; mem3[139]<=0; mem4[139]<=0;
mem1[140]<=0;  mem2[140]<=0; mem3[140]<=0; mem4[140]<=0;
mem1[141]<=0;  mem2[141]<=0; mem3[141]<=0; mem4[141]<=0;
mem1[142]<=0;  mem2[142]<=0; mem3[142]<=0; mem4[142]<=0;
mem1[143]<=0;  mem2[143]<=0; mem3[143]<=0; mem4[143]<=0;
mem1[144]<=0;  mem2[144]<=0; mem3[144]<=0; mem4[144]<=0;
mem1[145]<=0;  mem2[145]<=0; mem3[145]<=0; mem4[145]<=0;
mem1[146]<=0;  mem2[146]<=0; mem3[146]<=0; mem4[146]<=0;
mem1[147]<=0;  mem2[147]<=0; mem3[147]<=0; mem4[147]<=0;
mem1[148]<=0;  mem2[148]<=0; mem3[148]<=0; mem4[148]<=0;
mem1[149]<=0;  mem2[149]<=0; mem3[149]<=0; mem4[149]<=0;
mem1[150]<=0;  mem2[150]<=0; mem3[150]<=0; mem4[150]<=0;
mem1[151]<=0;  mem2[151]<=0; mem3[151]<=0; mem4[151]<=0;
mem1[152]<=0;  mem2[152]<=0; mem3[152]<=0; mem4[152]<=0;
mem1[153]<=0;  mem2[153]<=0; mem3[153]<=0; mem4[153]<=0;
mem1[154]<=0;  mem2[154]<=0; mem3[154]<=0; mem4[154]<=0;
mem1[155]<=0;  mem2[155]<=0; mem3[155]<=0; mem4[155]<=0;
mem1[156]<=0;  mem2[156]<=0; mem3[156]<=0; mem4[156]<=0;
mem1[157]<=0;  mem2[157]<=0; mem3[157]<=0; mem4[157]<=0;
mem1[158]<=0;  mem2[158]<=0; mem3[158]<=0; mem4[158]<=0;
mem1[159]<=0;  mem2[159]<=0; mem3[159]<=0; mem4[159]<=0;
mem1[160]<=0;  mem2[160]<=0; mem3[160]<=0; mem4[160]<=0;
mem1[161]<=0;  mem2[161]<=0; mem3[161]<=0; mem4[161]<=0;
mem1[162]<=0;  mem2[162]<=0; mem3[162]<=0; mem4[162]<=0;
mem1[163]<=0;  mem2[163]<=0; mem3[163]<=0; mem4[163]<=0;
mem1[164]<=0;  mem2[164]<=0; mem3[164]<=0; mem4[164]<=0;
mem1[165]<=0;  mem2[165]<=0; mem3[165]<=0; mem4[165]<=0;
mem1[166]<=0;  mem2[166]<=0; mem3[166]<=0; mem4[166]<=0;
mem1[167]<=0;  mem2[167]<=0; mem3[167]<=0; mem4[167]<=0;
mem1[168]<=0;  mem2[168]<=0; mem3[168]<=0; mem4[168]<=0;
mem1[169]<=0;  mem2[169]<=0; mem3[169]<=0; mem4[169]<=0;
mem1[170]<=0;  mem2[170]<=0; mem3[170]<=0; mem4[170]<=0;
mem1[171]<=0;  mem2[171]<=0; mem3[171]<=0; mem4[171]<=0;
mem1[172]<=0;  mem2[172]<=0; mem3[172]<=0; mem4[172]<=0;
mem1[173]<=0;  mem2[173]<=0; mem3[173]<=0; mem4[173]<=0;
mem1[174]<=0;  mem2[174]<=0; mem3[174]<=0; mem4[174]<=0;
mem1[175]<=0;  mem2[175]<=0; mem3[175]<=0; mem4[175]<=0;
mem1[176]<=0;  mem2[176]<=0; mem3[176]<=0; mem4[176]<=0;
mem1[177]<=0;  mem2[177]<=0; mem3[177]<=0; mem4[177]<=0;
mem1[178]<=0;  mem2[178]<=0; mem3[178]<=0; mem4[178]<=0;
mem1[179]<=0;  mem2[179]<=0; mem3[179]<=0; mem4[179]<=0;
mem1[180]<=0;  mem2[180]<=0; mem3[180]<=0; mem4[180]<=0;
mem1[181]<=0;  mem2[181]<=0; mem3[181]<=0; mem4[181]<=0;
mem1[182]<=0;  mem2[182]<=0; mem3[182]<=0; mem4[182]<=0;
mem1[183]<=0;  mem2[183]<=0; mem3[183]<=0; mem4[183]<=0;
mem1[184]<=0;  mem2[184]<=0; mem3[184]<=0; mem4[184]<=0;
mem1[185]<=0;  mem2[185]<=0; mem3[185]<=0; mem4[185]<=0;
mem1[186]<=0;  mem2[186]<=0; mem3[186]<=0; mem4[186]<=0;
mem1[187]<=0;  mem2[187]<=0; mem3[187]<=0; mem4[187]<=0;
mem1[188]<=0;  mem2[188]<=0; mem3[188]<=0; mem4[188]<=0;
mem1[189]<=0;  mem2[189]<=0; mem3[189]<=0; mem4[189]<=0;
mem1[190]<=0;  mem2[190]<=0; mem3[190]<=0; mem4[190]<=0;
mem1[191]<=0;  mem2[191]<=0; mem3[191]<=0; mem4[191]<=0;
mem1[192]<=0;  mem2[192]<=0; mem3[192]<=0; mem4[192]<=0;
mem1[193]<=0;  mem2[193]<=0; mem3[193]<=0; mem4[193]<=0;
mem1[194]<=0;  mem2[194]<=0; mem3[194]<=0; mem4[194]<=0;
mem1[195]<=0;  mem2[195]<=0; mem3[195]<=0; mem4[195]<=0;
mem1[196]<=0;  mem2[196]<=0; mem3[196]<=0; mem4[196]<=0;
mem1[197]<=0;  mem2[197]<=0; mem3[197]<=0; mem4[197]<=0;
mem1[198]<=0;  mem2[198]<=0; mem3[198]<=0; mem4[198]<=0;
mem1[199]<=0;  mem2[199]<=0; mem3[199]<=0; mem4[199]<=0;
mem1[200]<=0;  mem2[200]<=0; mem3[200]<=0; mem4[200]<=0;
mem1[201]<=0;  mem2[201]<=0; mem3[201]<=0; mem4[201]<=0;
mem1[202]<=0;  mem2[202]<=0; mem3[202]<=0; mem4[202]<=0;
mem1[203]<=0;  mem2[203]<=0; mem3[203]<=0; mem4[203]<=0;
mem1[204]<=0;  mem2[204]<=0; mem3[204]<=0; mem4[204]<=0;
mem1[205]<=0;  mem2[205]<=0; mem3[205]<=0; mem4[205]<=0;
mem1[206]<=0;  mem2[206]<=0; mem3[206]<=0; mem4[206]<=0;
mem1[207]<=0;  mem2[207]<=0; mem3[207]<=0; mem4[207]<=0;
mem1[208]<=0;  mem2[208]<=0; mem3[208]<=0; mem4[208]<=0;
mem1[209]<=0;  mem2[209]<=0; mem3[209]<=0; mem4[209]<=0;
mem1[210]<=0;  mem2[210]<=0; mem3[210]<=0; mem4[210]<=0;
mem1[211]<=0;  mem2[211]<=0; mem3[211]<=0; mem4[211]<=0;
mem1[212]<=0;  mem2[212]<=0; mem3[212]<=0; mem4[212]<=0;
mem1[213]<=0;  mem2[213]<=0; mem3[213]<=0; mem4[213]<=0;
mem1[214]<=0;  mem2[214]<=0; mem3[214]<=0; mem4[214]<=0;
mem1[215]<=0;  mem2[215]<=0; mem3[215]<=0; mem4[215]<=0;
mem1[216]<=0;  mem2[216]<=0; mem3[216]<=0; mem4[216]<=0;
mem1[217]<=0;  mem2[217]<=0; mem3[217]<=0; mem4[217]<=0;
mem1[218]<=0;  mem2[218]<=0; mem3[218]<=0; mem4[218]<=0;
mem1[219]<=0;  mem2[219]<=0; mem3[219]<=0; mem4[219]<=0;
mem1[220]<=0;  mem2[220]<=0; mem3[220]<=0; mem4[220]<=0;
mem1[221]<=0;  mem2[221]<=0; mem3[221]<=0; mem4[221]<=0;
mem1[222]<=0;  mem2[222]<=0; mem3[222]<=0; mem4[222]<=0;
mem1[223]<=0;  mem2[223]<=0; mem3[223]<=0; mem4[223]<=0;
mem1[224]<=0;  mem2[224]<=0; mem3[224]<=0; mem4[224]<=0;
mem1[225]<=0;  mem2[225]<=0; mem3[225]<=0; mem4[225]<=0;
mem1[226]<=0;  mem2[226]<=0; mem3[226]<=0; mem4[226]<=0;
mem1[227]<=0;  mem2[227]<=0; mem3[227]<=0; mem4[227]<=0;
mem1[228]<=0;  mem2[228]<=0; mem3[228]<=0; mem4[228]<=0;
mem1[229]<=0;  mem2[229]<=0; mem3[229]<=0; mem4[229]<=0;
mem1[230]<=0;  mem2[230]<=0; mem3[230]<=0; mem4[230]<=0;
mem1[231]<=0;  mem2[231]<=0; mem3[231]<=0; mem4[231]<=0;
mem1[232]<=0;  mem2[232]<=0; mem3[232]<=0; mem4[232]<=0;
mem1[233]<=0;  mem2[233]<=0; mem3[233]<=0; mem4[233]<=0;
mem1[234]<=0;  mem2[234]<=0; mem3[234]<=0; mem4[234]<=0;
mem1[235]<=0;  mem2[235]<=0; mem3[235]<=0; mem4[235]<=0;
mem1[236]<=0;  mem2[236]<=0; mem3[236]<=0; mem4[236]<=0;
mem1[237]<=0;  mem2[237]<=0; mem3[237]<=0; mem4[237]<=0;
mem1[238]<=0;  mem2[238]<=0; mem3[238]<=0; mem4[238]<=0;
mem1[239]<=0;  mem2[239]<=0; mem3[239]<=0; mem4[239]<=0;
mem1[240]<=0;  mem2[240]<=0; mem3[240]<=0; mem4[240]<=0;
mem1[241]<=0;  mem2[241]<=0; mem3[241]<=0; mem4[241]<=0;
mem1[242]<=0;  mem2[242]<=0; mem3[242]<=0; mem4[242]<=0;
mem1[243]<=0;  mem2[243]<=0; mem3[243]<=0; mem4[243]<=0;
mem1[244]<=0;  mem2[244]<=0; mem3[244]<=0; mem4[244]<=0;
mem1[245]<=0;  mem2[245]<=0; mem3[245]<=0; mem4[245]<=0;
mem1[246]<=0;  mem2[246]<=0; mem3[246]<=0; mem4[246]<=0;
mem1[247]<=0;  mem2[247]<=0; mem3[247]<=0; mem4[247]<=0;
mem1[248]<=0;  mem2[248]<=0; mem3[248]<=0; mem4[248]<=0;
mem1[249]<=0;  mem2[249]<=0; mem3[249]<=0; mem4[249]<=0;
mem1[250]<=0;  mem2[250]<=0; mem3[250]<=0; mem4[250]<=0;
mem1[251]<=0;  mem2[251]<=0; mem3[251]<=0; mem4[251]<=0;
mem1[252]<=0;  mem2[252]<=0; mem3[252]<=0; mem4[252]<=0;
mem1[253]<=0;  mem2[253]<=0; mem3[253]<=0; mem4[253]<=0;
mem1[254]<=0;  mem2[254]<=0; mem3[254]<=0; mem4[254]<=0;
mem1[255]<=0;  mem2[255]<=0; mem3[255]<=0; mem4[255]<=0;
mem1[256]<=0;  mem2[256]<=0; mem3[256]<=0; mem4[256]<=0;
mem1[257]<=0;  mem2[257]<=0; mem3[257]<=0; mem4[257]<=0;
mem1[258]<=0;  mem2[258]<=0; mem3[258]<=0; mem4[258]<=0;
mem1[259]<=0;  mem2[259]<=0; mem3[259]<=0; mem4[259]<=0;
mem1[260]<=0;  mem2[260]<=0; mem3[260]<=0; mem4[260]<=0;
mem1[261]<=0;  mem2[261]<=0; mem3[261]<=0; mem4[261]<=0;
mem1[262]<=0;  mem2[262]<=0; mem3[262]<=0; mem4[262]<=0;
mem1[263]<=0;  mem2[263]<=0; mem3[263]<=0; mem4[263]<=0;
mem1[264]<=0;  mem2[264]<=0; mem3[264]<=0; mem4[264]<=0;
mem1[265]<=0;  mem2[265]<=0; mem3[265]<=0; mem4[265]<=0;
mem1[266]<=0;  mem2[266]<=0; mem3[266]<=0; mem4[266]<=0;
mem1[267]<=0;  mem2[267]<=0; mem3[267]<=0; mem4[267]<=0;
mem1[268]<=0;  mem2[268]<=0; mem3[268]<=0; mem4[268]<=0;
mem1[269]<=0;  mem2[269]<=0; mem3[269]<=0; mem4[269]<=0;
mem1[270]<=0;  mem2[270]<=0; mem3[270]<=0; mem4[270]<=0;
mem1[271]<=0;  mem2[271]<=0; mem3[271]<=0; mem4[271]<=0;
mem1[272]<=0;  mem2[272]<=0; mem3[272]<=0; mem4[272]<=0;
mem1[273]<=0;  mem2[273]<=0; mem3[273]<=0; mem4[273]<=0;
mem1[274]<=0;  mem2[274]<=0; mem3[274]<=0; mem4[274]<=0;
mem1[275]<=0;  mem2[275]<=0; mem3[275]<=0; mem4[275]<=0;
mem1[276]<=0;  mem2[276]<=0; mem3[276]<=0; mem4[276]<=0;
mem1[277]<=0;  mem2[277]<=0; mem3[277]<=0; mem4[277]<=0;
mem1[278]<=0;  mem2[278]<=0; mem3[278]<=0; mem4[278]<=0;
mem1[279]<=0;  mem2[279]<=0; mem3[279]<=0; mem4[279]<=0;
mem1[280]<=0;  mem2[280]<=0; mem3[280]<=0; mem4[280]<=0;
mem1[281]<=0;  mem2[281]<=0; mem3[281]<=0; mem4[281]<=0;
mem1[282]<=0;  mem2[282]<=0; mem3[282]<=0; mem4[282]<=0;
mem1[283]<=0;  mem2[283]<=0; mem3[283]<=0; mem4[283]<=0;
mem1[284]<=0;  mem2[284]<=0; mem3[284]<=0; mem4[284]<=0;
mem1[285]<=0;  mem2[285]<=0; mem3[285]<=0; mem4[285]<=0;
mem1[286]<=0;  mem2[286]<=0; mem3[286]<=0; mem4[286]<=0;
mem1[287]<=0;  mem2[287]<=0; mem3[287]<=0; mem4[287]<=0;
mem1[288]<=0;  mem2[288]<=0; mem3[288]<=0; mem4[288]<=0;
mem1[289]<=0;  mem2[289]<=0; mem3[289]<=0; mem4[289]<=0;
mem1[290]<=0;  mem2[290]<=0; mem3[290]<=0; mem4[290]<=0;
mem1[291]<=0;  mem2[291]<=0; mem3[291]<=0; mem4[291]<=0;
mem1[292]<=0;  mem2[292]<=0; mem3[292]<=0; mem4[292]<=0;
mem1[293]<=0;  mem2[293]<=0; mem3[293]<=0; mem4[293]<=0;
mem1[294]<=0;  mem2[294]<=0; mem3[294]<=0; mem4[294]<=0;
mem1[295]<=0;  mem2[295]<=0; mem3[295]<=0; mem4[295]<=0;
mem1[296]<=0;  mem2[296]<=0; mem3[296]<=0; mem4[296]<=0;
mem1[297]<=0;  mem2[297]<=0; mem3[297]<=0; mem4[297]<=0;
mem1[298]<=0;  mem2[298]<=0; mem3[298]<=0; mem4[298]<=0;
mem1[299]<=0;  mem2[299]<=0; mem3[299]<=0; mem4[299]<=0;
mem1[300]<=0;  mem2[300]<=0; mem3[300]<=0; mem4[300]<=0;
mem1[301]<=0;  mem2[301]<=0; mem3[301]<=0; mem4[301]<=0;
mem1[302]<=0;  mem2[302]<=0; mem3[302]<=0; mem4[302]<=0;
mem1[303]<=0;  mem2[303]<=0; mem3[303]<=0; mem4[303]<=0;
mem1[304]<=0;  mem2[304]<=0; mem3[304]<=0; mem4[304]<=0;
mem1[305]<=0;  mem2[305]<=0; mem3[305]<=0; mem4[305]<=0;
mem1[306]<=0;  mem2[306]<=0; mem3[306]<=0; mem4[306]<=0;
mem1[307]<=0;  mem2[307]<=0; mem3[307]<=0; mem4[307]<=0;
mem1[308]<=0;  mem2[308]<=0; mem3[308]<=0; mem4[308]<=0;
mem1[309]<=0;  mem2[309]<=0; mem3[309]<=0; mem4[309]<=0;
mem1[310]<=0;  mem2[310]<=0; mem3[310]<=0; mem4[310]<=0;
mem1[311]<=0;  mem2[311]<=0; mem3[311]<=0; mem4[311]<=0;
mem1[312]<=0;  mem2[312]<=0; mem3[312]<=0; mem4[312]<=0;
mem1[313]<=0;  mem2[313]<=0; mem3[313]<=0; mem4[313]<=0;
mem1[314]<=0;  mem2[314]<=0; mem3[314]<=0; mem4[314]<=0;
mem1[315]<=0;  mem2[315]<=0; mem3[315]<=0; mem4[315]<=0;
mem1[316]<=0;  mem2[316]<=0; mem3[316]<=0; mem4[316]<=0;
mem1[317]<=0;  mem2[317]<=0; mem3[317]<=0; mem4[317]<=0;
mem1[318]<=0;  mem2[318]<=0; mem3[318]<=0; mem4[318]<=0;
mem1[319]<=0;  mem2[319]<=0; mem3[319]<=0; mem4[319]<=0;
mem1[320]<=0;  mem2[320]<=0; mem3[320]<=0; mem4[320]<=0;
mem1[321]<=0;  mem2[321]<=0; mem3[321]<=0; mem4[321]<=0;
mem1[322]<=0;  mem2[322]<=0; mem3[322]<=0; mem4[322]<=0;
mem1[323]<=0;  mem2[323]<=0; mem3[323]<=0; mem4[323]<=0;
mem1[324]<=0;  mem2[324]<=0; mem3[324]<=0; mem4[324]<=0;
mem1[325]<=0;  mem2[325]<=0; mem3[325]<=0; mem4[325]<=0;
mem1[326]<=0;  mem2[326]<=0; mem3[326]<=0; mem4[326]<=0;
mem1[327]<=0;  mem2[327]<=0; mem3[327]<=0; mem4[327]<=0;
mem1[328]<=0;  mem2[328]<=0; mem3[328]<=0; mem4[328]<=0;
mem1[329]<=0;  mem2[329]<=0; mem3[329]<=0; mem4[329]<=0;
mem1[330]<=0;  mem2[330]<=0; mem3[330]<=0; mem4[330]<=0;
mem1[331]<=0;  mem2[331]<=0; mem3[331]<=0; mem4[331]<=0;
mem1[332]<=0;  mem2[332]<=0; mem3[332]<=0; mem4[332]<=0;
mem1[333]<=0;  mem2[333]<=0; mem3[333]<=0; mem4[333]<=0;
mem1[334]<=0;  mem2[334]<=0; mem3[334]<=0; mem4[334]<=0;
mem1[335]<=0;  mem2[335]<=0; mem3[335]<=0; mem4[335]<=0;
mem1[336]<=0;  mem2[336]<=0; mem3[336]<=0; mem4[336]<=0;
mem1[337]<=0;  mem2[337]<=0; mem3[337]<=0; mem4[337]<=0;
mem1[338]<=0;  mem2[338]<=0; mem3[338]<=0; mem4[338]<=0;
mem1[339]<=0;  mem2[339]<=0; mem3[339]<=0; mem4[339]<=0;
mem1[340]<=0;  mem2[340]<=0; mem3[340]<=0; mem4[340]<=0;
mem1[341]<=0;  mem2[341]<=0; mem3[341]<=0; mem4[341]<=0;
mem1[342]<=0;  mem2[342]<=0; mem3[342]<=0; mem4[342]<=0;
mem1[343]<=0;  mem2[343]<=0; mem3[343]<=0; mem4[343]<=0;
mem1[344]<=0;  mem2[344]<=0; mem3[344]<=0; mem4[344]<=0;
mem1[345]<=0;  mem2[345]<=0; mem3[345]<=0; mem4[345]<=0;
mem1[346]<=0;  mem2[346]<=0; mem3[346]<=0; mem4[346]<=0;
mem1[347]<=0;  mem2[347]<=0; mem3[347]<=0; mem4[347]<=0;
mem1[348]<=0;  mem2[348]<=0; mem3[348]<=0; mem4[348]<=0;
mem1[349]<=0;  mem2[349]<=0; mem3[349]<=0; mem4[349]<=0;
mem1[350]<=0;  mem2[350]<=0; mem3[350]<=0; mem4[350]<=0;
mem1[351]<=0;  mem2[351]<=0; mem3[351]<=0; mem4[351]<=0;
mem1[352]<=0;  mem2[352]<=0; mem3[352]<=0; mem4[352]<=0;
mem1[353]<=0;  mem2[353]<=0; mem3[353]<=0; mem4[353]<=0;
mem1[354]<=0;  mem2[354]<=0; mem3[354]<=0; mem4[354]<=0;
mem1[355]<=0;  mem2[355]<=0; mem3[355]<=0; mem4[355]<=0;
mem1[356]<=0;  mem2[356]<=0; mem3[356]<=0; mem4[356]<=0;
mem1[357]<=0;  mem2[357]<=0; mem3[357]<=0; mem4[357]<=0;
mem1[358]<=0;  mem2[358]<=0; mem3[358]<=0; mem4[358]<=0;
mem1[359]<=0;  mem2[359]<=0; mem3[359]<=0; mem4[359]<=0;
mem1[360]<=0;  mem2[360]<=0; mem3[360]<=0; mem4[360]<=0;
mem1[361]<=0;  mem2[361]<=0; mem3[361]<=0; mem4[361]<=0;
mem1[362]<=0;  mem2[362]<=0; mem3[362]<=0; mem4[362]<=0;
mem1[363]<=0;  mem2[363]<=0; mem3[363]<=0; mem4[363]<=0;
mem1[364]<=0;  mem2[364]<=0; mem3[364]<=0; mem4[364]<=0;
mem1[365]<=0;  mem2[365]<=0; mem3[365]<=0; mem4[365]<=0;
mem1[366]<=0;  mem2[366]<=0; mem3[366]<=0; mem4[366]<=0;
mem1[367]<=0;  mem2[367]<=0; mem3[367]<=0; mem4[367]<=0;
mem1[368]<=0;  mem2[368]<=0; mem3[368]<=0; mem4[368]<=0;
mem1[369]<=0;  mem2[369]<=0; mem3[369]<=0; mem4[369]<=0;
mem1[370]<=0;  mem2[370]<=0; mem3[370]<=0; mem4[370]<=0;
mem1[371]<=0;  mem2[371]<=0; mem3[371]<=0; mem4[371]<=0;
mem1[372]<=0;  mem2[372]<=0; mem3[372]<=0; mem4[372]<=0;
mem1[373]<=0;  mem2[373]<=0; mem3[373]<=0; mem4[373]<=0;
mem1[374]<=0;  mem2[374]<=0; mem3[374]<=0; mem4[374]<=0;
mem1[375]<=0;  mem2[375]<=0; mem3[375]<=0; mem4[375]<=0;
mem1[376]<=0;  mem2[376]<=0; mem3[376]<=0; mem4[376]<=0;
mem1[377]<=0;  mem2[377]<=0; mem3[377]<=0; mem4[377]<=0;
mem1[378]<=0;  mem2[378]<=0; mem3[378]<=0; mem4[378]<=0;
mem1[379]<=0;  mem2[379]<=0; mem3[379]<=0; mem4[379]<=0;
mem1[380]<=0;  mem2[380]<=0; mem3[380]<=0; mem4[380]<=0;
mem1[381]<=0;  mem2[381]<=0; mem3[381]<=0; mem4[381]<=0;
mem1[382]<=0;  mem2[382]<=0; mem3[382]<=0; mem4[382]<=0;
mem1[383]<=0;  mem2[383]<=0; mem3[383]<=0; mem4[383]<=0;
mem1[384]<=0;  mem2[384]<=0; mem3[384]<=0; mem4[384]<=0;
mem1[385]<=0;  mem2[385]<=0; mem3[385]<=0; mem4[385]<=0;
mem1[386]<=0;  mem2[386]<=0; mem3[386]<=0; mem4[386]<=0;
mem1[387]<=0;  mem2[387]<=0; mem3[387]<=0; mem4[387]<=0;
mem1[388]<=0;  mem2[388]<=0; mem3[388]<=0; mem4[388]<=0;
mem1[389]<=0;  mem2[389]<=0; mem3[389]<=0; mem4[389]<=0;
mem1[390]<=0;  mem2[390]<=0; mem3[390]<=0; mem4[390]<=0;
mem1[391]<=0;  mem2[391]<=0; mem3[391]<=0; mem4[391]<=0;
mem1[392]<=0;  mem2[392]<=0; mem3[392]<=0; mem4[392]<=0;
mem1[393]<=0;  mem2[393]<=0; mem3[393]<=0; mem4[393]<=0;
mem1[394]<=0;  mem2[394]<=0; mem3[394]<=0; mem4[394]<=0;
mem1[395]<=0;  mem2[395]<=0; mem3[395]<=0; mem4[395]<=0;
mem1[396]<=0;  mem2[396]<=0; mem3[396]<=0; mem4[396]<=0;
mem1[397]<=0;  mem2[397]<=0; mem3[397]<=0; mem4[397]<=0;
mem1[398]<=0;  mem2[398]<=0; mem3[398]<=0; mem4[398]<=0;
mem1[399]<=0;  mem2[399]<=0; mem3[399]<=0; mem4[399]<=0;
mem1[400]<=0;  mem2[400]<=0; mem3[400]<=0; mem4[400]<=0;
mem1[401]<=0;  mem2[401]<=0; mem3[401]<=0; mem4[401]<=0;
mem1[402]<=0;  mem2[402]<=0; mem3[402]<=0; mem4[402]<=0;
mem1[403]<=0;  mem2[403]<=0; mem3[403]<=0; mem4[403]<=0;
mem1[404]<=0;  mem2[404]<=0; mem3[404]<=0; mem4[404]<=0;
mem1[405]<=0;  mem2[405]<=0; mem3[405]<=0; mem4[405]<=0;
mem1[406]<=0;  mem2[406]<=0; mem3[406]<=0; mem4[406]<=0;
mem1[407]<=0;  mem2[407]<=0; mem3[407]<=0; mem4[407]<=0;
mem1[408]<=0;  mem2[408]<=0; mem3[408]<=0; mem4[408]<=0;
mem1[409]<=0;  mem2[409]<=0; mem3[409]<=0; mem4[409]<=0;
mem1[410]<=0;  mem2[410]<=0; mem3[410]<=0; mem4[410]<=0;
mem1[411]<=0;  mem2[411]<=0; mem3[411]<=0; mem4[411]<=0;
mem1[412]<=0;  mem2[412]<=0; mem3[412]<=0; mem4[412]<=0;
mem1[413]<=0;  mem2[413]<=0; mem3[413]<=0; mem4[413]<=0;
mem1[414]<=0;  mem2[414]<=0; mem3[414]<=0; mem4[414]<=0;
mem1[415]<=0;  mem2[415]<=0; mem3[415]<=0; mem4[415]<=0;
mem1[416]<=0;  mem2[416]<=0; mem3[416]<=0; mem4[416]<=0;
mem1[417]<=0;  mem2[417]<=0; mem3[417]<=0; mem4[417]<=0;
mem1[418]<=0;  mem2[418]<=0; mem3[418]<=0; mem4[418]<=0;
mem1[419]<=0;  mem2[419]<=0; mem3[419]<=0; mem4[419]<=0;
mem1[420]<=0;  mem2[420]<=0; mem3[420]<=0; mem4[420]<=0;
mem1[421]<=0;  mem2[421]<=0; mem3[421]<=0; mem4[421]<=0;
mem1[422]<=0;  mem2[422]<=0; mem3[422]<=0; mem4[422]<=0;
mem1[423]<=0;  mem2[423]<=0; mem3[423]<=0; mem4[423]<=0;
mem1[424]<=0;  mem2[424]<=0; mem3[424]<=0; mem4[424]<=0;
mem1[425]<=0;  mem2[425]<=0; mem3[425]<=0; mem4[425]<=0;
mem1[426]<=0;  mem2[426]<=0; mem3[426]<=0; mem4[426]<=0;
mem1[427]<=0;  mem2[427]<=0; mem3[427]<=0; mem4[427]<=0;
mem1[428]<=0;  mem2[428]<=0; mem3[428]<=0; mem4[428]<=0;
mem1[429]<=0;  mem2[429]<=0; mem3[429]<=0; mem4[429]<=0;
mem1[430]<=0;  mem2[430]<=0; mem3[430]<=0; mem4[430]<=0;
mem1[431]<=0;  mem2[431]<=0; mem3[431]<=0; mem4[431]<=0;
mem1[432]<=0;  mem2[432]<=0; mem3[432]<=0; mem4[432]<=0;
mem1[433]<=0;  mem2[433]<=0; mem3[433]<=0; mem4[433]<=0;
mem1[434]<=0;  mem2[434]<=0; mem3[434]<=0; mem4[434]<=0;
mem1[435]<=0;  mem2[435]<=0; mem3[435]<=0; mem4[435]<=0;
mem1[436]<=0;  mem2[436]<=0; mem3[436]<=0; mem4[436]<=0;
mem1[437]<=0;  mem2[437]<=0; mem3[437]<=0; mem4[437]<=0;
mem1[438]<=0;  mem2[438]<=0; mem3[438]<=0; mem4[438]<=0;
mem1[439]<=0;  mem2[439]<=0; mem3[439]<=0; mem4[439]<=0;
mem1[440]<=0;  mem2[440]<=0; mem3[440]<=0; mem4[440]<=0;
mem1[441]<=0;  mem2[441]<=0; mem3[441]<=0; mem4[441]<=0;
mem1[442]<=0;  mem2[442]<=0; mem3[442]<=0; mem4[442]<=0;
mem1[443]<=0;  mem2[443]<=0; mem3[443]<=0; mem4[443]<=0;
mem1[444]<=0;  mem2[444]<=0; mem3[444]<=0; mem4[444]<=0;
mem1[445]<=0;  mem2[445]<=0; mem3[445]<=0; mem4[445]<=0;
mem1[446]<=0;  mem2[446]<=0; mem3[446]<=0; mem4[446]<=0;
mem1[447]<=0;  mem2[447]<=0; mem3[447]<=0; mem4[447]<=0;
mem1[448]<=0;  mem2[448]<=0; mem3[448]<=0; mem4[448]<=0;
mem1[449]<=0;  mem2[449]<=0; mem3[449]<=0; mem4[449]<=0;
mem1[450]<=0;  mem2[450]<=0; mem3[450]<=0; mem4[450]<=0;
mem1[451]<=0;  mem2[451]<=0; mem3[451]<=0; mem4[451]<=0;
mem1[452]<=0;  mem2[452]<=0; mem3[452]<=0; mem4[452]<=0;
mem1[453]<=0;  mem2[453]<=0; mem3[453]<=0; mem4[453]<=0;
mem1[454]<=0;  mem2[454]<=0; mem3[454]<=0; mem4[454]<=0;
mem1[455]<=0;  mem2[455]<=0; mem3[455]<=0; mem4[455]<=0;
mem1[456]<=0;  mem2[456]<=0; mem3[456]<=0; mem4[456]<=0;
mem1[457]<=0;  mem2[457]<=0; mem3[457]<=0; mem4[457]<=0;
mem1[458]<=0;  mem2[458]<=0; mem3[458]<=0; mem4[458]<=0;
mem1[459]<=0;  mem2[459]<=0; mem3[459]<=0; mem4[459]<=0;
mem1[460]<=0;  mem2[460]<=0; mem3[460]<=0; mem4[460]<=0;
mem1[461]<=0;  mem2[461]<=0; mem3[461]<=0; mem4[461]<=0;
mem1[462]<=0;  mem2[462]<=0; mem3[462]<=0; mem4[462]<=0;
mem1[463]<=0;  mem2[463]<=0; mem3[463]<=0; mem4[463]<=0;
mem1[464]<=0;  mem2[464]<=0; mem3[464]<=0; mem4[464]<=0;
mem1[465]<=0;  mem2[465]<=0; mem3[465]<=0; mem4[465]<=0;
mem1[466]<=0;  mem2[466]<=0; mem3[466]<=0; mem4[466]<=0;
mem1[467]<=0;  mem2[467]<=0; mem3[467]<=0; mem4[467]<=0;
mem1[468]<=0;  mem2[468]<=0; mem3[468]<=0; mem4[468]<=0;
mem1[469]<=0;  mem2[469]<=0; mem3[469]<=0; mem4[469]<=0;
mem1[470]<=0;  mem2[470]<=0; mem3[470]<=0; mem4[470]<=0;
mem1[471]<=0;  mem2[471]<=0; mem3[471]<=0; mem4[471]<=0;
mem1[472]<=0;  mem2[472]<=0; mem3[472]<=0; mem4[472]<=0;
mem1[473]<=0;  mem2[473]<=0; mem3[473]<=0; mem4[473]<=0;
mem1[474]<=0;  mem2[474]<=0; mem3[474]<=0; mem4[474]<=0;
mem1[475]<=0;  mem2[475]<=0; mem3[475]<=0; mem4[475]<=0;
mem1[476]<=0;  mem2[476]<=0; mem3[476]<=0; mem4[476]<=0;
mem1[477]<=0;  mem2[477]<=0; mem3[477]<=0; mem4[477]<=0;
mem1[478]<=0;  mem2[478]<=0; mem3[478]<=0; mem4[478]<=0;
mem1[479]<=0;  mem2[479]<=0; mem3[479]<=0; mem4[479]<=0;
mem1[480]<=0;  mem2[480]<=0; mem3[480]<=0; mem4[480]<=0;
mem1[481]<=0;  mem2[481]<=0; mem3[481]<=0; mem4[481]<=0;
mem1[482]<=0;  mem2[482]<=0; mem3[482]<=0; mem4[482]<=0;
mem1[483]<=0;  mem2[483]<=0; mem3[483]<=0; mem4[483]<=0;
mem1[484]<=0;  mem2[484]<=0; mem3[484]<=0; mem4[484]<=0;
mem1[485]<=0;  mem2[485]<=0; mem3[485]<=0; mem4[485]<=0;
mem1[486]<=0;  mem2[486]<=0; mem3[486]<=0; mem4[486]<=0;
mem1[487]<=0;  mem2[487]<=0; mem3[487]<=0; mem4[487]<=0;
mem1[488]<=0;  mem2[488]<=0; mem3[488]<=0; mem4[488]<=0;
mem1[489]<=0;  mem2[489]<=0; mem3[489]<=0; mem4[489]<=0;
mem1[490]<=0;  mem2[490]<=0; mem3[490]<=0; mem4[490]<=0;
mem1[491]<=0;  mem2[491]<=0; mem3[491]<=0; mem4[491]<=0;
mem1[492]<=0;  mem2[492]<=0; mem3[492]<=0; mem4[492]<=0;
mem1[493]<=0;  mem2[493]<=0; mem3[493]<=0; mem4[493]<=0;
mem1[494]<=0;  mem2[494]<=0; mem3[494]<=0; mem4[494]<=0;
mem1[495]<=0;  mem2[495]<=0; mem3[495]<=0; mem4[495]<=0;
mem1[496]<=0;  mem2[496]<=0; mem3[496]<=0; mem4[496]<=0;
mem1[497]<=0;  mem2[497]<=0; mem3[497]<=0; mem4[497]<=0;
mem1[498]<=0;  mem2[498]<=0; mem3[498]<=0; mem4[498]<=0;
mem1[499]<=0;  mem2[499]<=0; mem3[499]<=0; mem4[499]<=0;
mem1[500]<=0;  mem2[500]<=0; mem3[500]<=0; mem4[500]<=0;
mem1[501]<=0;  mem2[501]<=0; mem3[501]<=0; mem4[501]<=0;
mem1[502]<=0;  mem2[502]<=0; mem3[502]<=0; mem4[502]<=0;
mem1[503]<=0;  mem2[503]<=0; mem3[503]<=0; mem4[503]<=0;
mem1[504]<=0;  mem2[504]<=0; mem3[504]<=0; mem4[504]<=0;
mem1[505]<=0;  mem2[505]<=0; mem3[505]<=0; mem4[505]<=0;
mem1[506]<=0;  mem2[506]<=0; mem3[506]<=0; mem4[506]<=0;
mem1[507]<=0;  mem2[507]<=0; mem3[507]<=0; mem4[507]<=0;
mem1[508]<=0;  mem2[508]<=0; mem3[508]<=0; mem4[508]<=0;
mem1[509]<=0;  mem2[509]<=0; mem3[509]<=0; mem4[509]<=0;
mem1[510]<=0;  mem2[510]<=0; mem3[510]<=0; mem4[510]<=0;
mem1[511]<=0;  mem2[511]<=0; mem3[511]<=0; mem4[511]<=0;
mem1[512]<=0;  mem2[512]<=0; mem3[512]<=0; mem4[512]<=0;
mem1[513]<=0;  mem2[513]<=0; mem3[513]<=0; mem4[513]<=0;
mem1[514]<=0;  mem2[514]<=0; mem3[514]<=0; mem4[514]<=0;
mem1[515]<=0;  mem2[515]<=0; mem3[515]<=0; mem4[515]<=0;
mem1[516]<=0;  mem2[516]<=0; mem3[516]<=0; mem4[516]<=0;
mem1[517]<=0;  mem2[517]<=0; mem3[517]<=0; mem4[517]<=0;
mem1[518]<=0;  mem2[518]<=0; mem3[518]<=0; mem4[518]<=0;
mem1[519]<=0;  mem2[519]<=0; mem3[519]<=0; mem4[519]<=0;
mem1[520]<=0;  mem2[520]<=0; mem3[520]<=0; mem4[520]<=0;
mem1[521]<=0;  mem2[521]<=0; mem3[521]<=0; mem4[521]<=0;
mem1[522]<=0;  mem2[522]<=0; mem3[522]<=0; mem4[522]<=0;
mem1[523]<=0;  mem2[523]<=0; mem3[523]<=0; mem4[523]<=0;
mem1[524]<=0;  mem2[524]<=0; mem3[524]<=0; mem4[524]<=0;
mem1[525]<=0;  mem2[525]<=0; mem3[525]<=0; mem4[525]<=0;
mem1[526]<=0;  mem2[526]<=0; mem3[526]<=0; mem4[526]<=0;
mem1[527]<=0;  mem2[527]<=0; mem3[527]<=0; mem4[527]<=0;
mem1[528]<=0;  mem2[528]<=0; mem3[528]<=0; mem4[528]<=0;
mem1[529]<=0;  mem2[529]<=0; mem3[529]<=0; mem4[529]<=0;
mem1[530]<=0;  mem2[530]<=0; mem3[530]<=0; mem4[530]<=0;
mem1[531]<=0;  mem2[531]<=0; mem3[531]<=0; mem4[531]<=0;
mem1[532]<=0;  mem2[532]<=0; mem3[532]<=0; mem4[532]<=0;
mem1[533]<=0;  mem2[533]<=0; mem3[533]<=0; mem4[533]<=0;
mem1[534]<=0;  mem2[534]<=0; mem3[534]<=0; mem4[534]<=0;
mem1[535]<=0;  mem2[535]<=0; mem3[535]<=0; mem4[535]<=0;
mem1[536]<=0;  mem2[536]<=0; mem3[536]<=0; mem4[536]<=0;
mem1[537]<=0;  mem2[537]<=0; mem3[537]<=0; mem4[537]<=0;
mem1[538]<=0;  mem2[538]<=0; mem3[538]<=0; mem4[538]<=0;
mem1[539]<=0;  mem2[539]<=0; mem3[539]<=0; mem4[539]<=0;
mem1[540]<=0;  mem2[540]<=0; mem3[540]<=0; mem4[540]<=0;
mem1[541]<=0;  mem2[541]<=0; mem3[541]<=0; mem4[541]<=0;
mem1[542]<=0;  mem2[542]<=0; mem3[542]<=0; mem4[542]<=0;
mem1[543]<=0;  mem2[543]<=0; mem3[543]<=0; mem4[543]<=0;
mem1[544]<=0;  mem2[544]<=0; mem3[544]<=0; mem4[544]<=0;
mem1[545]<=0;  mem2[545]<=0; mem3[545]<=0; mem4[545]<=0;
mem1[546]<=0;  mem2[546]<=0; mem3[546]<=0; mem4[546]<=0;
mem1[547]<=0;  mem2[547]<=0; mem3[547]<=0; mem4[547]<=0;
mem1[548]<=0;  mem2[548]<=0; mem3[548]<=0; mem4[548]<=0;
mem1[549]<=0;  mem2[549]<=0; mem3[549]<=0; mem4[549]<=0;
mem1[550]<=0;  mem2[550]<=0; mem3[550]<=0; mem4[550]<=0;
mem1[551]<=0;  mem2[551]<=0; mem3[551]<=0; mem4[551]<=0;
mem1[552]<=0;  mem2[552]<=0; mem3[552]<=0; mem4[552]<=0;
mem1[553]<=0;  mem2[553]<=0; mem3[553]<=0; mem4[553]<=0;
mem1[554]<=0;  mem2[554]<=0; mem3[554]<=0; mem4[554]<=0;
mem1[555]<=0;  mem2[555]<=0; mem3[555]<=0; mem4[555]<=0;
mem1[556]<=0;  mem2[556]<=0; mem3[556]<=0; mem4[556]<=0;
mem1[557]<=0;  mem2[557]<=0; mem3[557]<=0; mem4[557]<=0;
mem1[558]<=0;  mem2[558]<=0; mem3[558]<=0; mem4[558]<=0;
mem1[559]<=0;  mem2[559]<=0; mem3[559]<=0; mem4[559]<=0;
mem1[560]<=0;  mem2[560]<=0; mem3[560]<=0; mem4[560]<=0;
mem1[561]<=0;  mem2[561]<=0; mem3[561]<=0; mem4[561]<=0;
mem1[562]<=0;  mem2[562]<=0; mem3[562]<=0; mem4[562]<=0;
mem1[563]<=0;  mem2[563]<=0; mem3[563]<=0; mem4[563]<=0;
mem1[564]<=0;  mem2[564]<=0; mem3[564]<=0; mem4[564]<=0;
mem1[565]<=0;  mem2[565]<=0; mem3[565]<=0; mem4[565]<=0;
mem1[566]<=0;  mem2[566]<=0; mem3[566]<=0; mem4[566]<=0;
mem1[567]<=0;  mem2[567]<=0; mem3[567]<=0; mem4[567]<=0;
mem1[568]<=0;  mem2[568]<=0; mem3[568]<=0; mem4[568]<=0;
mem1[569]<=0;  mem2[569]<=0; mem3[569]<=0; mem4[569]<=0;
mem1[570]<=0;  mem2[570]<=0; mem3[570]<=0; mem4[570]<=0;
mem1[571]<=0;  mem2[571]<=0; mem3[571]<=0; mem4[571]<=0;
mem1[572]<=0;  mem2[572]<=0; mem3[572]<=0; mem4[572]<=0;
mem1[573]<=0;  mem2[573]<=0; mem3[573]<=0; mem4[573]<=0;
mem1[574]<=0;  mem2[574]<=0; mem3[574]<=0; mem4[574]<=0;
mem1[575]<=0;  mem2[575]<=0; mem3[575]<=0; mem4[575]<=0;
mem1[576]<=0;  mem2[576]<=0; mem3[576]<=0; mem4[576]<=0;
mem1[577]<=0;  mem2[577]<=0; mem3[577]<=0; mem4[577]<=0;
mem1[578]<=0;  mem2[578]<=0; mem3[578]<=0; mem4[578]<=0;
mem1[579]<=0;  mem2[579]<=0; mem3[579]<=0; mem4[579]<=0;
mem1[580]<=0;  mem2[580]<=0; mem3[580]<=0; mem4[580]<=0;
mem1[581]<=0;  mem2[581]<=0; mem3[581]<=0; mem4[581]<=0;
mem1[582]<=0;  mem2[582]<=0; mem3[582]<=0; mem4[582]<=0;
mem1[583]<=0;  mem2[583]<=0; mem3[583]<=0; mem4[583]<=0;
mem1[584]<=0;  mem2[584]<=0; mem3[584]<=0; mem4[584]<=0;
mem1[585]<=0;  mem2[585]<=0; mem3[585]<=0; mem4[585]<=0;
mem1[586]<=0;  mem2[586]<=0; mem3[586]<=0; mem4[586]<=0;
mem1[587]<=0;  mem2[587]<=0; mem3[587]<=0; mem4[587]<=0;
mem1[588]<=0;  mem2[588]<=0; mem3[588]<=0; mem4[588]<=0;
mem1[589]<=0;  mem2[589]<=0; mem3[589]<=0; mem4[589]<=0;
mem1[590]<=0;  mem2[590]<=0; mem3[590]<=0; mem4[590]<=0;
mem1[591]<=0;  mem2[591]<=0; mem3[591]<=0; mem4[591]<=0;
mem1[592]<=0;  mem2[592]<=0; mem3[592]<=0; mem4[592]<=0;
mem1[593]<=0;  mem2[593]<=0; mem3[593]<=0; mem4[593]<=0;
mem1[594]<=0;  mem2[594]<=0; mem3[594]<=0; mem4[594]<=0;
mem1[595]<=0;  mem2[595]<=0; mem3[595]<=0; mem4[595]<=0;
mem1[596]<=0;  mem2[596]<=0; mem3[596]<=0; mem4[596]<=0;
mem1[597]<=0;  mem2[597]<=0; mem3[597]<=0; mem4[597]<=0;
mem1[598]<=0;  mem2[598]<=0; mem3[598]<=0; mem4[598]<=0;
mem1[599]<=0;  mem2[599]<=0; mem3[599]<=0; mem4[599]<=0;
mem1[600]<=0;  mem2[600]<=0; mem3[600]<=0; mem4[600]<=0;
mem1[601]<=0;  mem2[601]<=0; mem3[601]<=0; mem4[601]<=0;
mem1[602]<=0;  mem2[602]<=0; mem3[602]<=0; mem4[602]<=0;
mem1[603]<=0;  mem2[603]<=0; mem3[603]<=0; mem4[603]<=0;
mem1[604]<=0;  mem2[604]<=0; mem3[604]<=0; mem4[604]<=0;
mem1[605]<=0;  mem2[605]<=0; mem3[605]<=0; mem4[605]<=0;
mem1[606]<=0;  mem2[606]<=0; mem3[606]<=0; mem4[606]<=0;
mem1[607]<=0;  mem2[607]<=0; mem3[607]<=0; mem4[607]<=0;
mem1[608]<=0;  mem2[608]<=0; mem3[608]<=0; mem4[608]<=0;
mem1[609]<=0;  mem2[609]<=0; mem3[609]<=0; mem4[609]<=0;
mem1[610]<=0;  mem2[610]<=0; mem3[610]<=0; mem4[610]<=0;
mem1[611]<=0;  mem2[611]<=0; mem3[611]<=0; mem4[611]<=0;
mem1[612]<=0;  mem2[612]<=0; mem3[612]<=0; mem4[612]<=0;
mem1[613]<=0;  mem2[613]<=0; mem3[613]<=0; mem4[613]<=0;
mem1[614]<=0;  mem2[614]<=0; mem3[614]<=0; mem4[614]<=0;
mem1[615]<=0;  mem2[615]<=0; mem3[615]<=0; mem4[615]<=0;
mem1[616]<=0;  mem2[616]<=0; mem3[616]<=0; mem4[616]<=0;
mem1[617]<=0;  mem2[617]<=0; mem3[617]<=0; mem4[617]<=0;
mem1[618]<=0;  mem2[618]<=0; mem3[618]<=0; mem4[618]<=0;
mem1[619]<=0;  mem2[619]<=0; mem3[619]<=0; mem4[619]<=0;
mem1[620]<=0;  mem2[620]<=0; mem3[620]<=0; mem4[620]<=0;
mem1[621]<=0;  mem2[621]<=0; mem3[621]<=0; mem4[621]<=0;
mem1[622]<=0;  mem2[622]<=0; mem3[622]<=0; mem4[622]<=0;
mem1[623]<=0;  mem2[623]<=0; mem3[623]<=0; mem4[623]<=0;
mem1[624]<=0;  mem2[624]<=0; mem3[624]<=0; mem4[624]<=0;
mem1[625]<=0;  mem2[625]<=0; mem3[625]<=0; mem4[625]<=0;
mem1[626]<=0;  mem2[626]<=0; mem3[626]<=0; mem4[626]<=0;
mem1[627]<=0;  mem2[627]<=0; mem3[627]<=0; mem4[627]<=0;
mem1[628]<=0;  mem2[628]<=0; mem3[628]<=0; mem4[628]<=0;
mem1[629]<=0;  mem2[629]<=0; mem3[629]<=0; mem4[629]<=0;
mem1[630]<=0;  mem2[630]<=0; mem3[630]<=0; mem4[630]<=0;
mem1[631]<=0;  mem2[631]<=0; mem3[631]<=0; mem4[631]<=0;
mem1[632]<=0;  mem2[632]<=0; mem3[632]<=0; mem4[632]<=0;
mem1[633]<=0;  mem2[633]<=0; mem3[633]<=0; mem4[633]<=0;
mem1[634]<=0;  mem2[634]<=0; mem3[634]<=0; mem4[634]<=0;
mem1[635]<=0;  mem2[635]<=0; mem3[635]<=0; mem4[635]<=0;
mem1[636]<=0;  mem2[636]<=0; mem3[636]<=0; mem4[636]<=0;
mem1[637]<=0;  mem2[637]<=0; mem3[637]<=0; mem4[637]<=0;
mem1[638]<=0;  mem2[638]<=0; mem3[638]<=0; mem4[638]<=0;
mem1[639]<=0;  mem2[639]<=0; mem3[639]<=0; mem4[639]<=0;
mem1[640]<=0;  mem2[640]<=0; mem3[640]<=0; mem4[640]<=0;
mem1[641]<=0;  mem2[641]<=0; mem3[641]<=0; mem4[641]<=0;
mem1[642]<=0;  mem2[642]<=0; mem3[642]<=0; mem4[642]<=0;
mem1[643]<=0;  mem2[643]<=0; mem3[643]<=0; mem4[643]<=0;
mem1[644]<=0;  mem2[644]<=0; mem3[644]<=0; mem4[644]<=0;
mem1[645]<=0;  mem2[645]<=0; mem3[645]<=0; mem4[645]<=0;
mem1[646]<=0;  mem2[646]<=0; mem3[646]<=0; mem4[646]<=0;
mem1[647]<=0;  mem2[647]<=0; mem3[647]<=0; mem4[647]<=0;
mem1[648]<=0;  mem2[648]<=0; mem3[648]<=0; mem4[648]<=0;
mem1[649]<=0;  mem2[649]<=0; mem3[649]<=0; mem4[649]<=0;
mem1[650]<=0;  mem2[650]<=0; mem3[650]<=0; mem4[650]<=0;
mem1[651]<=0;  mem2[651]<=0; mem3[651]<=0; mem4[651]<=0;
mem1[652]<=0;  mem2[652]<=0; mem3[652]<=0; mem4[652]<=0;
mem1[653]<=0;  mem2[653]<=0; mem3[653]<=0; mem4[653]<=0;
mem1[654]<=0;  mem2[654]<=0; mem3[654]<=0; mem4[654]<=0;
mem1[655]<=0;  mem2[655]<=0; mem3[655]<=0; mem4[655]<=0;
mem1[656]<=0;  mem2[656]<=0; mem3[656]<=0; mem4[656]<=0;
mem1[657]<=0;  mem2[657]<=0; mem3[657]<=0; mem4[657]<=0;
mem1[658]<=0;  mem2[658]<=0; mem3[658]<=0; mem4[658]<=0;
mem1[659]<=0;  mem2[659]<=0; mem3[659]<=0; mem4[659]<=0;
mem1[660]<=0;  mem2[660]<=0; mem3[660]<=0; mem4[660]<=0;
mem1[661]<=0;  mem2[661]<=0; mem3[661]<=0; mem4[661]<=0;
mem1[662]<=0;  mem2[662]<=0; mem3[662]<=0; mem4[662]<=0;
mem1[663]<=0;  mem2[663]<=0; mem3[663]<=0; mem4[663]<=0;
mem1[664]<=0;  mem2[664]<=0; mem3[664]<=0; mem4[664]<=0;
mem1[665]<=0;  mem2[665]<=0; mem3[665]<=0; mem4[665]<=0;
mem1[666]<=0;  mem2[666]<=0; mem3[666]<=0; mem4[666]<=0;
mem1[667]<=0;  mem2[667]<=0; mem3[667]<=0; mem4[667]<=0;
mem1[668]<=0;  mem2[668]<=0; mem3[668]<=0; mem4[668]<=0;
mem1[669]<=0;  mem2[669]<=0; mem3[669]<=0; mem4[669]<=0;
mem1[670]<=0;  mem2[670]<=0; mem3[670]<=0; mem4[670]<=0;
mem1[671]<=0;  mem2[671]<=0; mem3[671]<=0; mem4[671]<=0;
mem1[672]<=0;  mem2[672]<=0; mem3[672]<=0; mem4[672]<=0;
mem1[673]<=0;  mem2[673]<=0; mem3[673]<=0; mem4[673]<=0;
mem1[674]<=0;  mem2[674]<=0; mem3[674]<=0; mem4[674]<=0;
mem1[675]<=0;  mem2[675]<=0; mem3[675]<=0; mem4[675]<=0;
mem1[676]<=0;  mem2[676]<=0; mem3[676]<=0; mem4[676]<=0;
mem1[677]<=0;  mem2[677]<=0; mem3[677]<=0; mem4[677]<=0;
mem1[678]<=0;  mem2[678]<=0; mem3[678]<=0; mem4[678]<=0;
mem1[679]<=0;  mem2[679]<=0; mem3[679]<=0; mem4[679]<=0;
mem1[680]<=0;  mem2[680]<=0; mem3[680]<=0; mem4[680]<=0;
mem1[681]<=0;  mem2[681]<=0; mem3[681]<=0; mem4[681]<=0;
mem1[682]<=0;  mem2[682]<=0; mem3[682]<=0; mem4[682]<=0;
mem1[683]<=0;  mem2[683]<=0; mem3[683]<=0; mem4[683]<=0;
mem1[684]<=0;  mem2[684]<=0; mem3[684]<=0; mem4[684]<=0;
mem1[685]<=0;  mem2[685]<=0; mem3[685]<=0; mem4[685]<=0;
mem1[686]<=0;  mem2[686]<=0; mem3[686]<=0; mem4[686]<=0;
mem1[687]<=0;  mem2[687]<=0; mem3[687]<=0; mem4[687]<=0;
mem1[688]<=0;  mem2[688]<=0; mem3[688]<=0; mem4[688]<=0;
mem1[689]<=0;  mem2[689]<=0; mem3[689]<=0; mem4[689]<=0;
mem1[690]<=0;  mem2[690]<=0; mem3[690]<=0; mem4[690]<=0;
mem1[691]<=0;  mem2[691]<=0; mem3[691]<=0; mem4[691]<=0;
mem1[692]<=0;  mem2[692]<=0; mem3[692]<=0; mem4[692]<=0;
mem1[693]<=0;  mem2[693]<=0; mem3[693]<=0; mem4[693]<=0;
mem1[694]<=0;  mem2[694]<=0; mem3[694]<=0; mem4[694]<=0;
mem1[695]<=0;  mem2[695]<=0; mem3[695]<=0; mem4[695]<=0;
mem1[696]<=0;  mem2[696]<=0; mem3[696]<=0; mem4[696]<=0;
mem1[697]<=0;  mem2[697]<=0; mem3[697]<=0; mem4[697]<=0;
mem1[698]<=0;  mem2[698]<=0; mem3[698]<=0; mem4[698]<=0;
mem1[699]<=0;  mem2[699]<=0; mem3[699]<=0; mem4[699]<=0;
mem1[700]<=0;  mem2[700]<=0; mem3[700]<=0; mem4[700]<=0;
mem1[701]<=0;  mem2[701]<=0; mem3[701]<=0; mem4[701]<=0;
mem1[702]<=0;  mem2[702]<=0; mem3[702]<=0; mem4[702]<=0;
mem1[703]<=0;  mem2[703]<=0; mem3[703]<=0; mem4[703]<=0;
mem1[704]<=0;  mem2[704]<=0; mem3[704]<=0; mem4[704]<=0;
mem1[705]<=0;  mem2[705]<=0; mem3[705]<=0; mem4[705]<=0;
mem1[706]<=0;  mem2[706]<=0; mem3[706]<=0; mem4[706]<=0;
mem1[707]<=0;  mem2[707]<=0; mem3[707]<=0; mem4[707]<=0;
mem1[708]<=0;  mem2[708]<=0; mem3[708]<=0; mem4[708]<=0;
mem1[709]<=0;  mem2[709]<=0; mem3[709]<=0; mem4[709]<=0;
mem1[710]<=0;  mem2[710]<=0; mem3[710]<=0; mem4[710]<=0;
mem1[711]<=0;  mem2[711]<=0; mem3[711]<=0; mem4[711]<=0;
mem1[712]<=0;  mem2[712]<=0; mem3[712]<=0; mem4[712]<=0;
mem1[713]<=0;  mem2[713]<=0; mem3[713]<=0; mem4[713]<=0;
mem1[714]<=0;  mem2[714]<=0; mem3[714]<=0; mem4[714]<=0;
mem1[715]<=0;  mem2[715]<=0; mem3[715]<=0; mem4[715]<=0;
mem1[716]<=0;  mem2[716]<=0; mem3[716]<=0; mem4[716]<=0;
mem1[717]<=0;  mem2[717]<=0; mem3[717]<=0; mem4[717]<=0;
mem1[718]<=0;  mem2[718]<=0; mem3[718]<=0; mem4[718]<=0;
mem1[719]<=0;  mem2[719]<=0; mem3[719]<=0; mem4[719]<=0;
mem1[720]<=0;  mem2[720]<=0; mem3[720]<=0; mem4[720]<=0;
mem1[721]<=0;  mem2[721]<=0; mem3[721]<=0; mem4[721]<=0;
mem1[722]<=0;  mem2[722]<=0; mem3[722]<=0; mem4[722]<=0;
mem1[723]<=0;  mem2[723]<=0; mem3[723]<=0; mem4[723]<=0;
mem1[724]<=0;  mem2[724]<=0; mem3[724]<=0; mem4[724]<=0;
mem1[725]<=0;  mem2[725]<=0; mem3[725]<=0; mem4[725]<=0;
mem1[726]<=0;  mem2[726]<=0; mem3[726]<=0; mem4[726]<=0;
mem1[727]<=0;  mem2[727]<=0; mem3[727]<=0; mem4[727]<=0;
mem1[728]<=0;  mem2[728]<=0; mem3[728]<=0; mem4[728]<=0;
mem1[729]<=0;  mem2[729]<=0; mem3[729]<=0; mem4[729]<=0;
mem1[730]<=0;  mem2[730]<=0; mem3[730]<=0; mem4[730]<=0;
mem1[731]<=0;  mem2[731]<=0; mem3[731]<=0; mem4[731]<=0;
mem1[732]<=0;  mem2[732]<=0; mem3[732]<=0; mem4[732]<=0;
mem1[733]<=0;  mem2[733]<=0; mem3[733]<=0; mem4[733]<=0;
mem1[734]<=0;  mem2[734]<=0; mem3[734]<=0; mem4[734]<=0;
mem1[735]<=0;  mem2[735]<=0; mem3[735]<=0; mem4[735]<=0;
mem1[736]<=0;  mem2[736]<=0; mem3[736]<=0; mem4[736]<=0;
mem1[737]<=0;  mem2[737]<=0; mem3[737]<=0; mem4[737]<=0;
mem1[738]<=0;  mem2[738]<=0; mem3[738]<=0; mem4[738]<=0;
mem1[739]<=0;  mem2[739]<=0; mem3[739]<=0; mem4[739]<=0;
mem1[740]<=0;  mem2[740]<=0; mem3[740]<=0; mem4[740]<=0;
mem1[741]<=0;  mem2[741]<=0; mem3[741]<=0; mem4[741]<=0;
mem1[742]<=0;  mem2[742]<=0; mem3[742]<=0; mem4[742]<=0;
mem1[743]<=0;  mem2[743]<=0; mem3[743]<=0; mem4[743]<=0;
mem1[744]<=0;  mem2[744]<=0; mem3[744]<=0; mem4[744]<=0;
mem1[745]<=0;  mem2[745]<=0; mem3[745]<=0; mem4[745]<=0;
mem1[746]<=0;  mem2[746]<=0; mem3[746]<=0; mem4[746]<=0;
mem1[747]<=0;  mem2[747]<=0; mem3[747]<=0; mem4[747]<=0;
mem1[748]<=0;  mem2[748]<=0; mem3[748]<=0; mem4[748]<=0;
mem1[749]<=0;  mem2[749]<=0; mem3[749]<=0; mem4[749]<=0;
mem1[750]<=0;  mem2[750]<=0; mem3[750]<=0; mem4[750]<=0;
mem1[751]<=0;  mem2[751]<=0; mem3[751]<=0; mem4[751]<=0;
mem1[752]<=0;  mem2[752]<=0; mem3[752]<=0; mem4[752]<=0;
mem1[753]<=0;  mem2[753]<=0; mem3[753]<=0; mem4[753]<=0;
mem1[754]<=0;  mem2[754]<=0; mem3[754]<=0; mem4[754]<=0;
mem1[755]<=0;  mem2[755]<=0; mem3[755]<=0; mem4[755]<=0;
mem1[756]<=0;  mem2[756]<=0; mem3[756]<=0; mem4[756]<=0;
mem1[757]<=0;  mem2[757]<=0; mem3[757]<=0; mem4[757]<=0;
mem1[758]<=0;  mem2[758]<=0; mem3[758]<=0; mem4[758]<=0;
mem1[759]<=0;  mem2[759]<=0; mem3[759]<=0; mem4[759]<=0;
mem1[760]<=0;  mem2[760]<=0; mem3[760]<=0; mem4[760]<=0;
mem1[761]<=0;  mem2[761]<=0; mem3[761]<=0; mem4[761]<=0;
mem1[762]<=0;  mem2[762]<=0; mem3[762]<=0; mem4[762]<=0;
mem1[763]<=0;  mem2[763]<=0; mem3[763]<=0; mem4[763]<=0;
mem1[764]<=0;  mem2[764]<=0; mem3[764]<=0; mem4[764]<=0;
mem1[765]<=0;  mem2[765]<=0; mem3[765]<=0; mem4[765]<=0;
mem1[766]<=0;  mem2[766]<=0; mem3[766]<=0; mem4[766]<=0;
mem1[767]<=0;  mem2[767]<=0; mem3[767]<=0; mem4[767]<=0;
mem1[768]<=0;  mem2[768]<=0; mem3[768]<=0; mem4[768]<=0;
mem1[769]<=0;  mem2[769]<=0; mem3[769]<=0; mem4[769]<=0;
mem1[770]<=0;  mem2[770]<=0; mem3[770]<=0; mem4[770]<=0;
mem1[771]<=0;  mem2[771]<=0; mem3[771]<=0; mem4[771]<=0;
mem1[772]<=0;  mem2[772]<=0; mem3[772]<=0; mem4[772]<=0;
mem1[773]<=0;  mem2[773]<=0; mem3[773]<=0; mem4[773]<=0;
mem1[774]<=0;  mem2[774]<=0; mem3[774]<=0; mem4[774]<=0;
mem1[775]<=0;  mem2[775]<=0; mem3[775]<=0; mem4[775]<=0;
mem1[776]<=0;  mem2[776]<=0; mem3[776]<=0; mem4[776]<=0;
mem1[777]<=0;  mem2[777]<=0; mem3[777]<=0; mem4[777]<=0;
mem1[778]<=0;  mem2[778]<=0; mem3[778]<=0; mem4[778]<=0;
mem1[779]<=0;  mem2[779]<=0; mem3[779]<=0; mem4[779]<=0;
mem1[780]<=0;  mem2[780]<=0; mem3[780]<=0; mem4[780]<=0;
mem1[781]<=0;  mem2[781]<=0; mem3[781]<=0; mem4[781]<=0;
mem1[782]<=0;  mem2[782]<=0; mem3[782]<=0; mem4[782]<=0;
mem1[783]<=0;  mem2[783]<=0; mem3[783]<=0; mem4[783]<=0;
mem1[784]<=0;  mem2[784]<=0; mem3[784]<=0; mem4[784]<=0;
mem1[785]<=0;  mem2[785]<=0; mem3[785]<=0; mem4[785]<=0;
mem1[786]<=0;  mem2[786]<=0; mem3[786]<=0; mem4[786]<=0;
mem1[787]<=0;  mem2[787]<=0; mem3[787]<=0; mem4[787]<=0;
mem1[788]<=0;  mem2[788]<=0; mem3[788]<=0; mem4[788]<=0;
mem1[789]<=0;  mem2[789]<=0; mem3[789]<=0; mem4[789]<=0;
mem1[790]<=0;  mem2[790]<=0; mem3[790]<=0; mem4[790]<=0;
mem1[791]<=0;  mem2[791]<=0; mem3[791]<=0; mem4[791]<=0;
mem1[792]<=0;  mem2[792]<=0; mem3[792]<=0; mem4[792]<=0;
mem1[793]<=0;  mem2[793]<=0; mem3[793]<=0; mem4[793]<=0;
mem1[794]<=0;  mem2[794]<=0; mem3[794]<=0; mem4[794]<=0;
mem1[795]<=0;  mem2[795]<=0; mem3[795]<=0; mem4[795]<=0;
mem1[796]<=0;  mem2[796]<=0; mem3[796]<=0; mem4[796]<=0;
mem1[797]<=0;  mem2[797]<=0; mem3[797]<=0; mem4[797]<=0;
mem1[798]<=0;  mem2[798]<=0; mem3[798]<=0; mem4[798]<=0;
mem1[799]<=0;  mem2[799]<=0; mem3[799]<=0; mem4[799]<=0;
mem1[800]<=0;  mem2[800]<=0; mem3[800]<=0; mem4[800]<=0;
mem1[801]<=0;  mem2[801]<=0; mem3[801]<=0; mem4[801]<=0;
mem1[802]<=0;  mem2[802]<=0; mem3[802]<=0; mem4[802]<=0;
mem1[803]<=0;  mem2[803]<=0; mem3[803]<=0; mem4[803]<=0;
mem1[804]<=0;  mem2[804]<=0; mem3[804]<=0; mem4[804]<=0;
mem1[805]<=0;  mem2[805]<=0; mem3[805]<=0; mem4[805]<=0;
mem1[806]<=0;  mem2[806]<=0; mem3[806]<=0; mem4[806]<=0;
mem1[807]<=0;  mem2[807]<=0; mem3[807]<=0; mem4[807]<=0;
mem1[808]<=0;  mem2[808]<=0; mem3[808]<=0; mem4[808]<=0;
mem1[809]<=0;  mem2[809]<=0; mem3[809]<=0; mem4[809]<=0;
mem1[810]<=0;  mem2[810]<=0; mem3[810]<=0; mem4[810]<=0;
mem1[811]<=0;  mem2[811]<=0; mem3[811]<=0; mem4[811]<=0;
mem1[812]<=0;  mem2[812]<=0; mem3[812]<=0; mem4[812]<=0;
mem1[813]<=0;  mem2[813]<=0; mem3[813]<=0; mem4[813]<=0;
mem1[814]<=0;  mem2[814]<=0; mem3[814]<=0; mem4[814]<=0;
mem1[815]<=0;  mem2[815]<=0; mem3[815]<=0; mem4[815]<=0;
mem1[816]<=0;  mem2[816]<=0; mem3[816]<=0; mem4[816]<=0;
mem1[817]<=0;  mem2[817]<=0; mem3[817]<=0; mem4[817]<=0;
mem1[818]<=0;  mem2[818]<=0; mem3[818]<=0; mem4[818]<=0;
mem1[819]<=0;  mem2[819]<=0; mem3[819]<=0; mem4[819]<=0;
mem1[820]<=0;  mem2[820]<=0; mem3[820]<=0; mem4[820]<=0;
mem1[821]<=0;  mem2[821]<=0; mem3[821]<=0; mem4[821]<=0;
mem1[822]<=0;  mem2[822]<=0; mem3[822]<=0; mem4[822]<=0;
mem1[823]<=0;  mem2[823]<=0; mem3[823]<=0; mem4[823]<=0;
mem1[824]<=0;  mem2[824]<=0; mem3[824]<=0; mem4[824]<=0;
mem1[825]<=0;  mem2[825]<=0; mem3[825]<=0; mem4[825]<=0;
mem1[826]<=0;  mem2[826]<=0; mem3[826]<=0; mem4[826]<=0;
mem1[827]<=0;  mem2[827]<=0; mem3[827]<=0; mem4[827]<=0;
mem1[828]<=0;  mem2[828]<=0; mem3[828]<=0; mem4[828]<=0;
mem1[829]<=0;  mem2[829]<=0; mem3[829]<=0; mem4[829]<=0;
mem1[830]<=0;  mem2[830]<=0; mem3[830]<=0; mem4[830]<=0;
mem1[831]<=0;  mem2[831]<=0; mem3[831]<=0; mem4[831]<=0;
mem1[832]<=0;  mem2[832]<=0; mem3[832]<=0; mem4[832]<=0;
mem1[833]<=0;  mem2[833]<=0; mem3[833]<=0; mem4[833]<=0;
mem1[834]<=0;  mem2[834]<=0; mem3[834]<=0; mem4[834]<=0;
mem1[835]<=0;  mem2[835]<=0; mem3[835]<=0; mem4[835]<=0;
mem1[836]<=0;  mem2[836]<=0; mem3[836]<=0; mem4[836]<=0;
mem1[837]<=0;  mem2[837]<=0; mem3[837]<=0; mem4[837]<=0;
mem1[838]<=0;  mem2[838]<=0; mem3[838]<=0; mem4[838]<=0;
mem1[839]<=0;  mem2[839]<=0; mem3[839]<=0; mem4[839]<=0;
mem1[840]<=0;  mem2[840]<=0; mem3[840]<=0; mem4[840]<=0;
mem1[841]<=0;  mem2[841]<=0; mem3[841]<=0; mem4[841]<=0;
mem1[842]<=0;  mem2[842]<=0; mem3[842]<=0; mem4[842]<=0;
mem1[843]<=0;  mem2[843]<=0; mem3[843]<=0; mem4[843]<=0;
mem1[844]<=0;  mem2[844]<=0; mem3[844]<=0; mem4[844]<=0;
mem1[845]<=0;  mem2[845]<=0; mem3[845]<=0; mem4[845]<=0;
mem1[846]<=0;  mem2[846]<=0; mem3[846]<=0; mem4[846]<=0;
mem1[847]<=0;  mem2[847]<=0; mem3[847]<=0; mem4[847]<=0;
mem1[848]<=0;  mem2[848]<=0; mem3[848]<=0; mem4[848]<=0;
mem1[849]<=0;  mem2[849]<=0; mem3[849]<=0; mem4[849]<=0;
mem1[850]<=0;  mem2[850]<=0; mem3[850]<=0; mem4[850]<=0;
mem1[851]<=0;  mem2[851]<=0; mem3[851]<=0; mem4[851]<=0;
mem1[852]<=0;  mem2[852]<=0; mem3[852]<=0; mem4[852]<=0;
mem1[853]<=0;  mem2[853]<=0; mem3[853]<=0; mem4[853]<=0;
mem1[854]<=0;  mem2[854]<=0; mem3[854]<=0; mem4[854]<=0;
mem1[855]<=0;  mem2[855]<=0; mem3[855]<=0; mem4[855]<=0;
mem1[856]<=0;  mem2[856]<=0; mem3[856]<=0; mem4[856]<=0;
mem1[857]<=0;  mem2[857]<=0; mem3[857]<=0; mem4[857]<=0;
mem1[858]<=0;  mem2[858]<=0; mem3[858]<=0; mem4[858]<=0;
mem1[859]<=0;  mem2[859]<=0; mem3[859]<=0; mem4[859]<=0;
mem1[860]<=0;  mem2[860]<=0; mem3[860]<=0; mem4[860]<=0;
mem1[861]<=0;  mem2[861]<=0; mem3[861]<=0; mem4[861]<=0;
mem1[862]<=0;  mem2[862]<=0; mem3[862]<=0; mem4[862]<=0;
mem1[863]<=0;  mem2[863]<=0; mem3[863]<=0; mem4[863]<=0;
mem1[864]<=0;  mem2[864]<=0; mem3[864]<=0; mem4[864]<=0;
mem1[865]<=0;  mem2[865]<=0; mem3[865]<=0; mem4[865]<=0;
mem1[866]<=0;  mem2[866]<=0; mem3[866]<=0; mem4[866]<=0;
mem1[867]<=0;  mem2[867]<=0; mem3[867]<=0; mem4[867]<=0;
mem1[868]<=0;  mem2[868]<=0; mem3[868]<=0; mem4[868]<=0;
mem1[869]<=0;  mem2[869]<=0; mem3[869]<=0; mem4[869]<=0;
mem1[870]<=0;  mem2[870]<=0; mem3[870]<=0; mem4[870]<=0;
mem1[871]<=0;  mem2[871]<=0; mem3[871]<=0; mem4[871]<=0;
mem1[872]<=0;  mem2[872]<=0; mem3[872]<=0; mem4[872]<=0;
mem1[873]<=0;  mem2[873]<=0; mem3[873]<=0; mem4[873]<=0;
mem1[874]<=0;  mem2[874]<=0; mem3[874]<=0; mem4[874]<=0;
mem1[875]<=0;  mem2[875]<=0; mem3[875]<=0; mem4[875]<=0;
mem1[876]<=0;  mem2[876]<=0; mem3[876]<=0; mem4[876]<=0;
mem1[877]<=0;  mem2[877]<=0; mem3[877]<=0; mem4[877]<=0;
mem1[878]<=0;  mem2[878]<=0; mem3[878]<=0; mem4[878]<=0;
mem1[879]<=0;  mem2[879]<=0; mem3[879]<=0; mem4[879]<=0;
mem1[880]<=0;  mem2[880]<=0; mem3[880]<=0; mem4[880]<=0;
mem1[881]<=0;  mem2[881]<=0; mem3[881]<=0; mem4[881]<=0;
mem1[882]<=0;  mem2[882]<=0; mem3[882]<=0; mem4[882]<=0;
mem1[883]<=0;  mem2[883]<=0; mem3[883]<=0; mem4[883]<=0;
mem1[884]<=0;  mem2[884]<=0; mem3[884]<=0; mem4[884]<=0;
mem1[885]<=0;  mem2[885]<=0; mem3[885]<=0; mem4[885]<=0;
mem1[886]<=0;  mem2[886]<=0; mem3[886]<=0; mem4[886]<=0;
mem1[887]<=0;  mem2[887]<=0; mem3[887]<=0; mem4[887]<=0;
mem1[888]<=0;  mem2[888]<=0; mem3[888]<=0; mem4[888]<=0;
mem1[889]<=0;  mem2[889]<=0; mem3[889]<=0; mem4[889]<=0;
mem1[890]<=0;  mem2[890]<=0; mem3[890]<=0; mem4[890]<=0;
mem1[891]<=0;  mem2[891]<=0; mem3[891]<=0; mem4[891]<=0;
mem1[892]<=0;  mem2[892]<=0; mem3[892]<=0; mem4[892]<=0;
mem1[893]<=0;  mem2[893]<=0; mem3[893]<=0; mem4[893]<=0;
mem1[894]<=0;  mem2[894]<=0; mem3[894]<=0; mem4[894]<=0;
mem1[895]<=0;  mem2[895]<=0; mem3[895]<=0; mem4[895]<=0;
mem1[896]<=0;  mem2[896]<=0; mem3[896]<=0; mem4[896]<=0;
mem1[897]<=0;  mem2[897]<=0; mem3[897]<=0; mem4[897]<=0;
mem1[898]<=0;  mem2[898]<=0; mem3[898]<=0; mem4[898]<=0;
mem1[899]<=0;  mem2[899]<=0; mem3[899]<=0; mem4[899]<=0;
mem1[900]<=0;  mem2[900]<=0; mem3[900]<=0; mem4[900]<=0;
mem1[901]<=0;  mem2[901]<=0; mem3[901]<=0; mem4[901]<=0;
mem1[902]<=0;  mem2[902]<=0; mem3[902]<=0; mem4[902]<=0;
mem1[903]<=0;  mem2[903]<=0; mem3[903]<=0; mem4[903]<=0;
mem1[904]<=0;  mem2[904]<=0; mem3[904]<=0; mem4[904]<=0;
mem1[905]<=0;  mem2[905]<=0; mem3[905]<=0; mem4[905]<=0;
mem1[906]<=0;  mem2[906]<=0; mem3[906]<=0; mem4[906]<=0;
mem1[907]<=0;  mem2[907]<=0; mem3[907]<=0; mem4[907]<=0;
mem1[908]<=0;  mem2[908]<=0; mem3[908]<=0; mem4[908]<=0;
mem1[909]<=0;  mem2[909]<=0; mem3[909]<=0; mem4[909]<=0;
mem1[910]<=0;  mem2[910]<=0; mem3[910]<=0; mem4[910]<=0;
mem1[911]<=0;  mem2[911]<=0; mem3[911]<=0; mem4[911]<=0;
mem1[912]<=0;  mem2[912]<=0; mem3[912]<=0; mem4[912]<=0;
mem1[913]<=0;  mem2[913]<=0; mem3[913]<=0; mem4[913]<=0;
mem1[914]<=0;  mem2[914]<=0; mem3[914]<=0; mem4[914]<=0;
mem1[915]<=0;  mem2[915]<=0; mem3[915]<=0; mem4[915]<=0;
mem1[916]<=0;  mem2[916]<=0; mem3[916]<=0; mem4[916]<=0;
mem1[917]<=0;  mem2[917]<=0; mem3[917]<=0; mem4[917]<=0;
mem1[918]<=0;  mem2[918]<=0; mem3[918]<=0; mem4[918]<=0;
mem1[919]<=0;  mem2[919]<=0; mem3[919]<=0; mem4[919]<=0;
mem1[920]<=0;  mem2[920]<=0; mem3[920]<=0; mem4[920]<=0;
mem1[921]<=0;  mem2[921]<=0; mem3[921]<=0; mem4[921]<=0;
mem1[922]<=0;  mem2[922]<=0; mem3[922]<=0; mem4[922]<=0;
mem1[923]<=0;  mem2[923]<=0; mem3[923]<=0; mem4[923]<=0;
mem1[924]<=0;  mem2[924]<=0; mem3[924]<=0; mem4[924]<=0;
mem1[925]<=0;  mem2[925]<=0; mem3[925]<=0; mem4[925]<=0;
mem1[926]<=0;  mem2[926]<=0; mem3[926]<=0; mem4[926]<=0;
mem1[927]<=0;  mem2[927]<=0; mem3[927]<=0; mem4[927]<=0;
mem1[928]<=0;  mem2[928]<=0; mem3[928]<=0; mem4[928]<=0;
mem1[929]<=0;  mem2[929]<=0; mem3[929]<=0; mem4[929]<=0;
mem1[930]<=0;  mem2[930]<=0; mem3[930]<=0; mem4[930]<=0;
mem1[931]<=0;  mem2[931]<=0; mem3[931]<=0; mem4[931]<=0;
mem1[932]<=0;  mem2[932]<=0; mem3[932]<=0; mem4[932]<=0;
mem1[933]<=0;  mem2[933]<=0; mem3[933]<=0; mem4[933]<=0;
mem1[934]<=0;  mem2[934]<=0; mem3[934]<=0; mem4[934]<=0;
mem1[935]<=0;  mem2[935]<=0; mem3[935]<=0; mem4[935]<=0;
mem1[936]<=0;  mem2[936]<=0; mem3[936]<=0; mem4[936]<=0;
mem1[937]<=0;  mem2[937]<=0; mem3[937]<=0; mem4[937]<=0;
mem1[938]<=0;  mem2[938]<=0; mem3[938]<=0; mem4[938]<=0;
mem1[939]<=0;  mem2[939]<=0; mem3[939]<=0; mem4[939]<=0;
mem1[940]<=0;  mem2[940]<=0; mem3[940]<=0; mem4[940]<=0;
mem1[941]<=0;  mem2[941]<=0; mem3[941]<=0; mem4[941]<=0;
mem1[942]<=0;  mem2[942]<=0; mem3[942]<=0; mem4[942]<=0;
mem1[943]<=0;  mem2[943]<=0; mem3[943]<=0; mem4[943]<=0;
mem1[944]<=0;  mem2[944]<=0; mem3[944]<=0; mem4[944]<=0;
mem1[945]<=0;  mem2[945]<=0; mem3[945]<=0; mem4[945]<=0;
mem1[946]<=0;  mem2[946]<=0; mem3[946]<=0; mem4[946]<=0;
mem1[947]<=0;  mem2[947]<=0; mem3[947]<=0; mem4[947]<=0;
mem1[948]<=0;  mem2[948]<=0; mem3[948]<=0; mem4[948]<=0;
mem1[949]<=0;  mem2[949]<=0; mem3[949]<=0; mem4[949]<=0;
mem1[950]<=0;  mem2[950]<=0; mem3[950]<=0; mem4[950]<=0;
mem1[951]<=0;  mem2[951]<=0; mem3[951]<=0; mem4[951]<=0;
mem1[952]<=0;  mem2[952]<=0; mem3[952]<=0; mem4[952]<=0;
mem1[953]<=0;  mem2[953]<=0; mem3[953]<=0; mem4[953]<=0;
mem1[954]<=0;  mem2[954]<=0; mem3[954]<=0; mem4[954]<=0;
mem1[955]<=0;  mem2[955]<=0; mem3[955]<=0; mem4[955]<=0;
mem1[956]<=0;  mem2[956]<=0; mem3[956]<=0; mem4[956]<=0;
mem1[957]<=0;  mem2[957]<=0; mem3[957]<=0; mem4[957]<=0;
mem1[958]<=0;  mem2[958]<=0; mem3[958]<=0; mem4[958]<=0;
mem1[959]<=0;  mem2[959]<=0; mem3[959]<=0; mem4[959]<=0;
mem1[960]<=0;  mem2[960]<=0; mem3[960]<=0; mem4[960]<=0;
mem1[961]<=0;  mem2[961]<=0; mem3[961]<=0; mem4[961]<=0;
mem1[962]<=0;  mem2[962]<=0; mem3[962]<=0; mem4[962]<=0;
mem1[963]<=0;  mem2[963]<=0; mem3[963]<=0; mem4[963]<=0;
mem1[964]<=0;  mem2[964]<=0; mem3[964]<=0; mem4[964]<=0;
mem1[965]<=0;  mem2[965]<=0; mem3[965]<=0; mem4[965]<=0;
mem1[966]<=0;  mem2[966]<=0; mem3[966]<=0; mem4[966]<=0;
mem1[967]<=0;  mem2[967]<=0; mem3[967]<=0; mem4[967]<=0;
mem1[968]<=0;  mem2[968]<=0; mem3[968]<=0; mem4[968]<=0;
mem1[969]<=0;  mem2[969]<=0; mem3[969]<=0; mem4[969]<=0;
mem1[970]<=0;  mem2[970]<=0; mem3[970]<=0; mem4[970]<=0;
mem1[971]<=0;  mem2[971]<=0; mem3[971]<=0; mem4[971]<=0;
mem1[972]<=0;  mem2[972]<=0; mem3[972]<=0; mem4[972]<=0;
mem1[973]<=0;  mem2[973]<=0; mem3[973]<=0; mem4[973]<=0;
mem1[974]<=0;  mem2[974]<=0; mem3[974]<=0; mem4[974]<=0;
mem1[975]<=0;  mem2[975]<=0; mem3[975]<=0; mem4[975]<=0;
mem1[976]<=0;  mem2[976]<=0; mem3[976]<=0; mem4[976]<=0;
mem1[977]<=0;  mem2[977]<=0; mem3[977]<=0; mem4[977]<=0;
mem1[978]<=0;  mem2[978]<=0; mem3[978]<=0; mem4[978]<=0;
mem1[979]<=0;  mem2[979]<=0; mem3[979]<=0; mem4[979]<=0;
mem1[980]<=0;  mem2[980]<=0; mem3[980]<=0; mem4[980]<=0;
mem1[981]<=0;  mem2[981]<=0; mem3[981]<=0; mem4[981]<=0;
mem1[982]<=0;  mem2[982]<=0; mem3[982]<=0; mem4[982]<=0;
mem1[983]<=0;  mem2[983]<=0; mem3[983]<=0; mem4[983]<=0;
mem1[984]<=0;  mem2[984]<=0; mem3[984]<=0; mem4[984]<=0;
mem1[985]<=0;  mem2[985]<=0; mem3[985]<=0; mem4[985]<=0;
mem1[986]<=0;  mem2[986]<=0; mem3[986]<=0; mem4[986]<=0;
mem1[987]<=0;  mem2[987]<=0; mem3[987]<=0; mem4[987]<=0;
mem1[988]<=0;  mem2[988]<=0; mem3[988]<=0; mem4[988]<=0;
mem1[989]<=0;  mem2[989]<=0; mem3[989]<=0; mem4[989]<=0;
mem1[990]<=0;  mem2[990]<=0; mem3[990]<=0; mem4[990]<=0;
mem1[991]<=0;  mem2[991]<=0; mem3[991]<=0; mem4[991]<=0;
mem1[992]<=0;  mem2[992]<=0; mem3[992]<=0; mem4[992]<=0;
mem1[993]<=0;  mem2[993]<=0; mem3[993]<=0; mem4[993]<=0;
mem1[994]<=0;  mem2[994]<=0; mem3[994]<=0; mem4[994]<=0;
mem1[995]<=0;  mem2[995]<=0; mem3[995]<=0; mem4[995]<=0;
mem1[996]<=0;  mem2[996]<=0; mem3[996]<=0; mem4[996]<=0;
mem1[997]<=0;  mem2[997]<=0; mem3[997]<=0; mem4[997]<=0;
mem1[998]<=0;  mem2[998]<=0; mem3[998]<=0; mem4[998]<=0;
mem1[999]<=0;  mem2[999]<=0; mem3[999]<=0; mem4[999]<=0;
mem1[1000]<=0;  mem2[1000]<=0; mem3[1000]<=0; mem4[1000]<=0;
mem1[1001]<=0;  mem2[1001]<=0; mem3[1001]<=0; mem4[1001]<=0;
mem1[1002]<=0;  mem2[1002]<=0; mem3[1002]<=0; mem4[1002]<=0;
mem1[1003]<=0;  mem2[1003]<=0; mem3[1003]<=0; mem4[1003]<=0;
mem1[1004]<=0;  mem2[1004]<=0; mem3[1004]<=0; mem4[1004]<=0;
mem1[1005]<=0;  mem2[1005]<=0; mem3[1005]<=0; mem4[1005]<=0;
mem1[1006]<=0;  mem2[1006]<=0; mem3[1006]<=0; mem4[1006]<=0;
mem1[1007]<=0;  mem2[1007]<=0; mem3[1007]<=0; mem4[1007]<=0;
mem1[1008]<=0;  mem2[1008]<=0; mem3[1008]<=0; mem4[1008]<=0;
mem1[1009]<=0;  mem2[1009]<=0; mem3[1009]<=0; mem4[1009]<=0;
mem1[1010]<=0;  mem2[1010]<=0; mem3[1010]<=0; mem4[1010]<=0;
mem1[1011]<=0;  mem2[1011]<=0; mem3[1011]<=0; mem4[1011]<=0;
mem1[1012]<=0;  mem2[1012]<=0; mem3[1012]<=0; mem4[1012]<=0;
mem1[1013]<=0;  mem2[1013]<=0; mem3[1013]<=0; mem4[1013]<=0;
mem1[1014]<=0;  mem2[1014]<=0; mem3[1014]<=0; mem4[1014]<=0;
mem1[1015]<=0;  mem2[1015]<=0; mem3[1015]<=0; mem4[1015]<=0;
mem1[1016]<=0;  mem2[1016]<=0; mem3[1016]<=0; mem4[1016]<=0;
mem1[1017]<=0;  mem2[1017]<=0; mem3[1017]<=0; mem4[1017]<=0;
mem1[1018]<=0;  mem2[1018]<=0; mem3[1018]<=0; mem4[1018]<=0;
mem1[1019]<=0;  mem2[1019]<=0; mem3[1019]<=0; mem4[1019]<=0;
mem1[1020]<=0;  mem2[1020]<=0; mem3[1020]<=0; mem4[1020]<=0;
mem1[1021]<=0;  mem2[1021]<=0; mem3[1021]<=0; mem4[1021]<=0;
mem1[1022]<=0;  mem2[1022]<=0; mem3[1022]<=0; mem4[1022]<=0;
mem1[1023]<=0;  mem2[1023]<=0; mem3[1023]<=0; mem4[1023]<=0;
end

endmodule
